module Top_remcm_mini (
	ext_end_read, 
	ext_end_comp, 
	ext_end_send, 
	ext_enable, 
	ext_comp, 
	ext_send, 
	ext_kx, 
	ext_ky, 
	ext_W, 
	ext_H, 
	ext_xin, 
	ext_coe, 
	ext_psum1, 
	ext_psum2, 
	wen_coe_fifo, 
	coe_wfull, 
	wen_xin_fifo, 
	xin_wfull, 
	ren_psum_fifo, 
	psum_rempty, 
	ext_clk, 
	int_clk, 
	ext_rst_n, 
	int_rst_n, 
	VCCK, 
	GNDK);
   output ext_end_read;
   output ext_end_comp;
   output ext_end_send;
   input ext_enable;
   input ext_comp;
   input ext_send;
   input [1:0] ext_kx;
   input [1:0] ext_ky;
   input [3:0] ext_W;
   input [3:0] ext_H;
   input [7:0] ext_xin;
   input [7:0] ext_coe;
   output [20:0] ext_psum1;
   output [20:0] ext_psum2;
   input wen_coe_fifo;
   output coe_wfull;
   input wen_xin_fifo;
   output xin_wfull;
   input ren_psum_fifo;
   output psum_rempty;
   input ext_clk;
   input int_clk;
   input ext_rst_n;
   input int_rst_n;

   // Internal wires
   wire VSS;
   wire VDD;
   wire n3845;
   wire n3846;
   wire n3847;
   wire coe_rempty;
   wire xin_rempty;
   wire psum_wfull;
   wire wen_coe;
   wire wen_x;
   wire xen1;
   wire xen4;
   wire coen;
   wire adden;
   wire adden_sec;
   wire sel_ccp;
   wire int_end_read;
   wire int_end_comp;
   wire int_end_send;
   wire int_enable;
   wire int_comp;
   wire int_send;
   wire Mcntl_flag;
   wire Mcntl_Mcntldata_N453;
   wire Mcntl_Mcntldata_comp_psum;
   wire Msyncin_Msynkxy_0__synkx_sync2;
   wire Msyncin_Msynkxy_0__synkx_sync1;
   wire Mfifo_coe_M_ffmem_mem_15__0_;
   wire Mfifo_coe_M_ffmem_mem_15__1_;
   wire Mfifo_coe_M_ffmem_mem_15__2_;
   wire Mfifo_coe_M_ffmem_mem_15__3_;
   wire Mfifo_coe_M_ffmem_mem_15__4_;
   wire Mfifo_coe_M_ffmem_mem_15__5_;
   wire Mfifo_coe_M_ffmem_mem_15__6_;
   wire Mfifo_coe_M_ffmem_mem_15__7_;
   wire Mfifo_coe_M_ffmem_mem_14__0_;
   wire Mfifo_coe_M_ffmem_mem_14__1_;
   wire Mfifo_coe_M_ffmem_mem_14__2_;
   wire Mfifo_coe_M_ffmem_mem_14__3_;
   wire Mfifo_coe_M_ffmem_mem_14__4_;
   wire Mfifo_coe_M_ffmem_mem_14__5_;
   wire Mfifo_coe_M_ffmem_mem_14__6_;
   wire Mfifo_coe_M_ffmem_mem_14__7_;
   wire Mfifo_coe_M_ffmem_mem_13__0_;
   wire Mfifo_coe_M_ffmem_mem_13__1_;
   wire Mfifo_coe_M_ffmem_mem_13__2_;
   wire Mfifo_coe_M_ffmem_mem_13__3_;
   wire Mfifo_coe_M_ffmem_mem_13__4_;
   wire Mfifo_coe_M_ffmem_mem_13__5_;
   wire Mfifo_coe_M_ffmem_mem_13__6_;
   wire Mfifo_coe_M_ffmem_mem_13__7_;
   wire Mfifo_coe_M_ffmem_mem_12__0_;
   wire Mfifo_coe_M_ffmem_mem_12__1_;
   wire Mfifo_coe_M_ffmem_mem_12__2_;
   wire Mfifo_coe_M_ffmem_mem_12__3_;
   wire Mfifo_coe_M_ffmem_mem_12__4_;
   wire Mfifo_coe_M_ffmem_mem_12__5_;
   wire Mfifo_coe_M_ffmem_mem_12__6_;
   wire Mfifo_coe_M_ffmem_mem_12__7_;
   wire Mfifo_coe_M_ffmem_mem_11__0_;
   wire Mfifo_coe_M_ffmem_mem_11__1_;
   wire Mfifo_coe_M_ffmem_mem_11__2_;
   wire Mfifo_coe_M_ffmem_mem_11__3_;
   wire Mfifo_coe_M_ffmem_mem_11__4_;
   wire Mfifo_coe_M_ffmem_mem_11__5_;
   wire Mfifo_coe_M_ffmem_mem_11__6_;
   wire Mfifo_coe_M_ffmem_mem_11__7_;
   wire Mfifo_coe_M_ffmem_mem_10__0_;
   wire Mfifo_coe_M_ffmem_mem_10__1_;
   wire Mfifo_coe_M_ffmem_mem_10__2_;
   wire Mfifo_coe_M_ffmem_mem_10__3_;
   wire Mfifo_coe_M_ffmem_mem_10__4_;
   wire Mfifo_coe_M_ffmem_mem_10__5_;
   wire Mfifo_coe_M_ffmem_mem_10__6_;
   wire Mfifo_coe_M_ffmem_mem_10__7_;
   wire Mfifo_coe_M_ffmem_mem_9__0_;
   wire Mfifo_coe_M_ffmem_mem_9__1_;
   wire Mfifo_coe_M_ffmem_mem_9__2_;
   wire Mfifo_coe_M_ffmem_mem_9__3_;
   wire Mfifo_coe_M_ffmem_mem_9__4_;
   wire Mfifo_coe_M_ffmem_mem_9__5_;
   wire Mfifo_coe_M_ffmem_mem_9__6_;
   wire Mfifo_coe_M_ffmem_mem_9__7_;
   wire Mfifo_coe_M_ffmem_mem_8__0_;
   wire Mfifo_coe_M_ffmem_mem_8__1_;
   wire Mfifo_coe_M_ffmem_mem_8__2_;
   wire Mfifo_coe_M_ffmem_mem_8__3_;
   wire Mfifo_coe_M_ffmem_mem_8__4_;
   wire Mfifo_coe_M_ffmem_mem_8__5_;
   wire Mfifo_coe_M_ffmem_mem_8__6_;
   wire Mfifo_coe_M_ffmem_mem_8__7_;
   wire Mfifo_coe_M_ffmem_mem_7__0_;
   wire Mfifo_coe_M_ffmem_mem_7__1_;
   wire Mfifo_coe_M_ffmem_mem_7__2_;
   wire Mfifo_coe_M_ffmem_mem_7__3_;
   wire Mfifo_coe_M_ffmem_mem_7__4_;
   wire Mfifo_coe_M_ffmem_mem_7__5_;
   wire Mfifo_coe_M_ffmem_mem_7__6_;
   wire Mfifo_coe_M_ffmem_mem_7__7_;
   wire Mfifo_coe_M_ffmem_mem_6__0_;
   wire Mfifo_coe_M_ffmem_mem_6__1_;
   wire Mfifo_coe_M_ffmem_mem_6__2_;
   wire Mfifo_coe_M_ffmem_mem_6__3_;
   wire Mfifo_coe_M_ffmem_mem_6__4_;
   wire Mfifo_coe_M_ffmem_mem_6__5_;
   wire Mfifo_coe_M_ffmem_mem_6__6_;
   wire Mfifo_coe_M_ffmem_mem_6__7_;
   wire Mfifo_coe_M_ffmem_mem_5__0_;
   wire Mfifo_coe_M_ffmem_mem_5__1_;
   wire Mfifo_coe_M_ffmem_mem_5__2_;
   wire Mfifo_coe_M_ffmem_mem_5__3_;
   wire Mfifo_coe_M_ffmem_mem_5__4_;
   wire Mfifo_coe_M_ffmem_mem_5__5_;
   wire Mfifo_coe_M_ffmem_mem_5__6_;
   wire Mfifo_coe_M_ffmem_mem_5__7_;
   wire Mfifo_coe_M_ffmem_mem_4__0_;
   wire Mfifo_coe_M_ffmem_mem_4__1_;
   wire Mfifo_coe_M_ffmem_mem_4__2_;
   wire Mfifo_coe_M_ffmem_mem_4__3_;
   wire Mfifo_coe_M_ffmem_mem_4__4_;
   wire Mfifo_coe_M_ffmem_mem_4__5_;
   wire Mfifo_coe_M_ffmem_mem_4__6_;
   wire Mfifo_coe_M_ffmem_mem_4__7_;
   wire Mfifo_coe_M_ffmem_mem_3__0_;
   wire Mfifo_coe_M_ffmem_mem_3__1_;
   wire Mfifo_coe_M_ffmem_mem_3__2_;
   wire Mfifo_coe_M_ffmem_mem_3__3_;
   wire Mfifo_coe_M_ffmem_mem_3__4_;
   wire Mfifo_coe_M_ffmem_mem_3__5_;
   wire Mfifo_coe_M_ffmem_mem_3__6_;
   wire Mfifo_coe_M_ffmem_mem_3__7_;
   wire Mfifo_coe_M_ffmem_mem_2__0_;
   wire Mfifo_coe_M_ffmem_mem_2__1_;
   wire Mfifo_coe_M_ffmem_mem_2__2_;
   wire Mfifo_coe_M_ffmem_mem_2__3_;
   wire Mfifo_coe_M_ffmem_mem_2__4_;
   wire Mfifo_coe_M_ffmem_mem_2__5_;
   wire Mfifo_coe_M_ffmem_mem_2__6_;
   wire Mfifo_coe_M_ffmem_mem_2__7_;
   wire Mfifo_coe_M_ffmem_mem_1__0_;
   wire Mfifo_coe_M_ffmem_mem_1__1_;
   wire Mfifo_coe_M_ffmem_mem_1__2_;
   wire Mfifo_coe_M_ffmem_mem_1__3_;
   wire Mfifo_coe_M_ffmem_mem_1__4_;
   wire Mfifo_coe_M_ffmem_mem_1__5_;
   wire Mfifo_coe_M_ffmem_mem_1__6_;
   wire Mfifo_coe_M_ffmem_mem_1__7_;
   wire Mfifo_coe_M_ffmem_mem_0__0_;
   wire Mfifo_coe_M_ffmem_mem_0__1_;
   wire Mfifo_coe_M_ffmem_mem_0__2_;
   wire Mfifo_coe_M_ffmem_mem_0__3_;
   wire Mfifo_coe_M_ffmem_mem_0__4_;
   wire Mfifo_coe_M_ffmem_mem_0__5_;
   wire Mfifo_coe_M_ffmem_mem_0__6_;
   wire Mfifo_coe_M_ffmem_mem_0__7_;
   wire Mfifo_coe_M_rptr_rempty_val;
   wire Mfifo_coe_M_rptr_N1;
   wire Mfifo_coe_M_wptr_wfull_val;
   wire Mfifo_psum_M_ffmem_N117;
   wire Mfifo_psum_M_ffmem_N116;
   wire Mfifo_psum_M_ffmem_N115;
   wire Mfifo_psum_M_ffmem_N114;
   wire Mfifo_psum_M_ffmem_N113;
   wire Mfifo_psum_M_ffmem_N112;
   wire Mfifo_psum_M_ffmem_N111;
   wire Mfifo_psum_M_ffmem_N110;
   wire Mfifo_psum_M_ffmem_N109;
   wire Mfifo_psum_M_ffmem_N108;
   wire Mfifo_psum_M_ffmem_N107;
   wire Mfifo_psum_M_ffmem_N106;
   wire Mfifo_psum_M_ffmem_N105;
   wire Mfifo_psum_M_ffmem_N104;
   wire Mfifo_psum_M_ffmem_N103;
   wire Mfifo_psum_M_ffmem_N102;
   wire Mfifo_psum_M_ffmem_N101;
   wire Mfifo_psum_M_ffmem_N100;
   wire Mfifo_psum_M_ffmem_N99;
   wire Mfifo_psum_M_ffmem_N98;
   wire Mfifo_psum_M_ffmem_N97;
   wire Mfifo_psum_M_ffmem_N96;
   wire Mfifo_psum_M_ffmem_N95;
   wire Mfifo_psum_M_ffmem_N94;
   wire Mfifo_psum_M_ffmem_N93;
   wire Mfifo_psum_M_ffmem_N92;
   wire Mfifo_psum_M_ffmem_N91;
   wire Mfifo_psum_M_ffmem_N90;
   wire Mfifo_psum_M_ffmem_N89;
   wire Mfifo_psum_M_ffmem_N88;
   wire Mfifo_psum_M_ffmem_N87;
   wire Mfifo_psum_M_ffmem_N86;
   wire Mfifo_psum_M_ffmem_N85;
   wire Mfifo_psum_M_ffmem_N84;
   wire Mfifo_psum_M_ffmem_N83;
   wire Mfifo_psum_M_ffmem_N82;
   wire Mfifo_psum_M_ffmem_N81;
   wire Mfifo_psum_M_ffmem_N80;
   wire Mfifo_psum_M_ffmem_N79;
   wire Mfifo_psum_M_ffmem_N78;
   wire Mfifo_psum_M_ffmem_N77;
   wire Mfifo_psum_M_ffmem_N76;
   wire Mfifo_psum_M_ffmem_mem_15__0_;
   wire Mfifo_psum_M_ffmem_mem_15__1_;
   wire Mfifo_psum_M_ffmem_mem_15__2_;
   wire Mfifo_psum_M_ffmem_mem_15__3_;
   wire Mfifo_psum_M_ffmem_mem_15__4_;
   wire Mfifo_psum_M_ffmem_mem_15__5_;
   wire Mfifo_psum_M_ffmem_mem_15__6_;
   wire Mfifo_psum_M_ffmem_mem_15__7_;
   wire Mfifo_psum_M_ffmem_mem_15__8_;
   wire Mfifo_psum_M_ffmem_mem_15__9_;
   wire Mfifo_psum_M_ffmem_mem_15__10_;
   wire Mfifo_psum_M_ffmem_mem_15__11_;
   wire Mfifo_psum_M_ffmem_mem_15__12_;
   wire Mfifo_psum_M_ffmem_mem_15__13_;
   wire Mfifo_psum_M_ffmem_mem_15__14_;
   wire Mfifo_psum_M_ffmem_mem_15__15_;
   wire Mfifo_psum_M_ffmem_mem_15__16_;
   wire Mfifo_psum_M_ffmem_mem_15__17_;
   wire Mfifo_psum_M_ffmem_mem_15__18_;
   wire Mfifo_psum_M_ffmem_mem_15__19_;
   wire Mfifo_psum_M_ffmem_mem_15__20_;
   wire Mfifo_psum_M_ffmem_mem_15__21_;
   wire Mfifo_psum_M_ffmem_mem_15__22_;
   wire Mfifo_psum_M_ffmem_mem_15__23_;
   wire Mfifo_psum_M_ffmem_mem_15__24_;
   wire Mfifo_psum_M_ffmem_mem_15__25_;
   wire Mfifo_psum_M_ffmem_mem_15__26_;
   wire Mfifo_psum_M_ffmem_mem_15__27_;
   wire Mfifo_psum_M_ffmem_mem_15__28_;
   wire Mfifo_psum_M_ffmem_mem_15__29_;
   wire Mfifo_psum_M_ffmem_mem_15__30_;
   wire Mfifo_psum_M_ffmem_mem_15__31_;
   wire Mfifo_psum_M_ffmem_mem_15__32_;
   wire Mfifo_psum_M_ffmem_mem_15__33_;
   wire Mfifo_psum_M_ffmem_mem_15__34_;
   wire Mfifo_psum_M_ffmem_mem_15__35_;
   wire Mfifo_psum_M_ffmem_mem_15__36_;
   wire Mfifo_psum_M_ffmem_mem_15__37_;
   wire Mfifo_psum_M_ffmem_mem_15__38_;
   wire Mfifo_psum_M_ffmem_mem_15__39_;
   wire Mfifo_psum_M_ffmem_mem_15__40_;
   wire Mfifo_psum_M_ffmem_mem_15__41_;
   wire Mfifo_psum_M_ffmem_mem_14__0_;
   wire Mfifo_psum_M_ffmem_mem_14__1_;
   wire Mfifo_psum_M_ffmem_mem_14__2_;
   wire Mfifo_psum_M_ffmem_mem_14__3_;
   wire Mfifo_psum_M_ffmem_mem_14__4_;
   wire Mfifo_psum_M_ffmem_mem_14__5_;
   wire Mfifo_psum_M_ffmem_mem_14__6_;
   wire Mfifo_psum_M_ffmem_mem_14__7_;
   wire Mfifo_psum_M_ffmem_mem_14__8_;
   wire Mfifo_psum_M_ffmem_mem_14__9_;
   wire Mfifo_psum_M_ffmem_mem_14__10_;
   wire Mfifo_psum_M_ffmem_mem_14__11_;
   wire Mfifo_psum_M_ffmem_mem_14__12_;
   wire Mfifo_psum_M_ffmem_mem_14__13_;
   wire Mfifo_psum_M_ffmem_mem_14__14_;
   wire Mfifo_psum_M_ffmem_mem_14__15_;
   wire Mfifo_psum_M_ffmem_mem_14__16_;
   wire Mfifo_psum_M_ffmem_mem_14__17_;
   wire Mfifo_psum_M_ffmem_mem_14__18_;
   wire Mfifo_psum_M_ffmem_mem_14__19_;
   wire Mfifo_psum_M_ffmem_mem_14__20_;
   wire Mfifo_psum_M_ffmem_mem_14__21_;
   wire Mfifo_psum_M_ffmem_mem_14__22_;
   wire Mfifo_psum_M_ffmem_mem_14__23_;
   wire Mfifo_psum_M_ffmem_mem_14__24_;
   wire Mfifo_psum_M_ffmem_mem_14__25_;
   wire Mfifo_psum_M_ffmem_mem_14__26_;
   wire Mfifo_psum_M_ffmem_mem_14__27_;
   wire Mfifo_psum_M_ffmem_mem_14__28_;
   wire Mfifo_psum_M_ffmem_mem_14__29_;
   wire Mfifo_psum_M_ffmem_mem_14__30_;
   wire Mfifo_psum_M_ffmem_mem_14__31_;
   wire Mfifo_psum_M_ffmem_mem_14__32_;
   wire Mfifo_psum_M_ffmem_mem_14__33_;
   wire Mfifo_psum_M_ffmem_mem_14__34_;
   wire Mfifo_psum_M_ffmem_mem_14__35_;
   wire Mfifo_psum_M_ffmem_mem_14__36_;
   wire Mfifo_psum_M_ffmem_mem_14__37_;
   wire Mfifo_psum_M_ffmem_mem_14__38_;
   wire Mfifo_psum_M_ffmem_mem_14__39_;
   wire Mfifo_psum_M_ffmem_mem_14__40_;
   wire Mfifo_psum_M_ffmem_mem_14__41_;
   wire Mfifo_psum_M_ffmem_mem_13__0_;
   wire Mfifo_psum_M_ffmem_mem_13__1_;
   wire Mfifo_psum_M_ffmem_mem_13__2_;
   wire Mfifo_psum_M_ffmem_mem_13__3_;
   wire Mfifo_psum_M_ffmem_mem_13__4_;
   wire Mfifo_psum_M_ffmem_mem_13__5_;
   wire Mfifo_psum_M_ffmem_mem_13__6_;
   wire Mfifo_psum_M_ffmem_mem_13__7_;
   wire Mfifo_psum_M_ffmem_mem_13__8_;
   wire Mfifo_psum_M_ffmem_mem_13__9_;
   wire Mfifo_psum_M_ffmem_mem_13__10_;
   wire Mfifo_psum_M_ffmem_mem_13__11_;
   wire Mfifo_psum_M_ffmem_mem_13__12_;
   wire Mfifo_psum_M_ffmem_mem_13__13_;
   wire Mfifo_psum_M_ffmem_mem_13__14_;
   wire Mfifo_psum_M_ffmem_mem_13__15_;
   wire Mfifo_psum_M_ffmem_mem_13__16_;
   wire Mfifo_psum_M_ffmem_mem_13__17_;
   wire Mfifo_psum_M_ffmem_mem_13__18_;
   wire Mfifo_psum_M_ffmem_mem_13__19_;
   wire Mfifo_psum_M_ffmem_mem_13__20_;
   wire Mfifo_psum_M_ffmem_mem_13__21_;
   wire Mfifo_psum_M_ffmem_mem_13__22_;
   wire Mfifo_psum_M_ffmem_mem_13__23_;
   wire Mfifo_psum_M_ffmem_mem_13__24_;
   wire Mfifo_psum_M_ffmem_mem_13__25_;
   wire Mfifo_psum_M_ffmem_mem_13__26_;
   wire Mfifo_psum_M_ffmem_mem_13__27_;
   wire Mfifo_psum_M_ffmem_mem_13__28_;
   wire Mfifo_psum_M_ffmem_mem_13__29_;
   wire Mfifo_psum_M_ffmem_mem_13__30_;
   wire Mfifo_psum_M_ffmem_mem_13__31_;
   wire Mfifo_psum_M_ffmem_mem_13__32_;
   wire Mfifo_psum_M_ffmem_mem_13__33_;
   wire Mfifo_psum_M_ffmem_mem_13__34_;
   wire Mfifo_psum_M_ffmem_mem_13__35_;
   wire Mfifo_psum_M_ffmem_mem_13__36_;
   wire Mfifo_psum_M_ffmem_mem_13__37_;
   wire Mfifo_psum_M_ffmem_mem_13__38_;
   wire Mfifo_psum_M_ffmem_mem_13__39_;
   wire Mfifo_psum_M_ffmem_mem_13__40_;
   wire Mfifo_psum_M_ffmem_mem_13__41_;
   wire Mfifo_psum_M_ffmem_mem_12__0_;
   wire Mfifo_psum_M_ffmem_mem_12__1_;
   wire Mfifo_psum_M_ffmem_mem_12__2_;
   wire Mfifo_psum_M_ffmem_mem_12__3_;
   wire Mfifo_psum_M_ffmem_mem_12__4_;
   wire Mfifo_psum_M_ffmem_mem_12__5_;
   wire Mfifo_psum_M_ffmem_mem_12__6_;
   wire Mfifo_psum_M_ffmem_mem_12__7_;
   wire Mfifo_psum_M_ffmem_mem_12__8_;
   wire Mfifo_psum_M_ffmem_mem_12__9_;
   wire Mfifo_psum_M_ffmem_mem_12__10_;
   wire Mfifo_psum_M_ffmem_mem_12__11_;
   wire Mfifo_psum_M_ffmem_mem_12__12_;
   wire Mfifo_psum_M_ffmem_mem_12__13_;
   wire Mfifo_psum_M_ffmem_mem_12__14_;
   wire Mfifo_psum_M_ffmem_mem_12__15_;
   wire Mfifo_psum_M_ffmem_mem_12__16_;
   wire Mfifo_psum_M_ffmem_mem_12__17_;
   wire Mfifo_psum_M_ffmem_mem_12__18_;
   wire Mfifo_psum_M_ffmem_mem_12__19_;
   wire Mfifo_psum_M_ffmem_mem_12__20_;
   wire Mfifo_psum_M_ffmem_mem_12__21_;
   wire Mfifo_psum_M_ffmem_mem_12__22_;
   wire Mfifo_psum_M_ffmem_mem_12__23_;
   wire Mfifo_psum_M_ffmem_mem_12__24_;
   wire Mfifo_psum_M_ffmem_mem_12__25_;
   wire Mfifo_psum_M_ffmem_mem_12__26_;
   wire Mfifo_psum_M_ffmem_mem_12__27_;
   wire Mfifo_psum_M_ffmem_mem_12__28_;
   wire Mfifo_psum_M_ffmem_mem_12__29_;
   wire Mfifo_psum_M_ffmem_mem_12__30_;
   wire Mfifo_psum_M_ffmem_mem_12__31_;
   wire Mfifo_psum_M_ffmem_mem_12__32_;
   wire Mfifo_psum_M_ffmem_mem_12__33_;
   wire Mfifo_psum_M_ffmem_mem_12__34_;
   wire Mfifo_psum_M_ffmem_mem_12__35_;
   wire Mfifo_psum_M_ffmem_mem_12__36_;
   wire Mfifo_psum_M_ffmem_mem_12__37_;
   wire Mfifo_psum_M_ffmem_mem_12__38_;
   wire Mfifo_psum_M_ffmem_mem_12__39_;
   wire Mfifo_psum_M_ffmem_mem_12__40_;
   wire Mfifo_psum_M_ffmem_mem_12__41_;
   wire Mfifo_psum_M_ffmem_mem_11__0_;
   wire Mfifo_psum_M_ffmem_mem_11__1_;
   wire Mfifo_psum_M_ffmem_mem_11__2_;
   wire Mfifo_psum_M_ffmem_mem_11__3_;
   wire Mfifo_psum_M_ffmem_mem_11__4_;
   wire Mfifo_psum_M_ffmem_mem_11__5_;
   wire Mfifo_psum_M_ffmem_mem_11__6_;
   wire Mfifo_psum_M_ffmem_mem_11__7_;
   wire Mfifo_psum_M_ffmem_mem_11__8_;
   wire Mfifo_psum_M_ffmem_mem_11__9_;
   wire Mfifo_psum_M_ffmem_mem_11__10_;
   wire Mfifo_psum_M_ffmem_mem_11__11_;
   wire Mfifo_psum_M_ffmem_mem_11__12_;
   wire Mfifo_psum_M_ffmem_mem_11__13_;
   wire Mfifo_psum_M_ffmem_mem_11__14_;
   wire Mfifo_psum_M_ffmem_mem_11__15_;
   wire Mfifo_psum_M_ffmem_mem_11__16_;
   wire Mfifo_psum_M_ffmem_mem_11__17_;
   wire Mfifo_psum_M_ffmem_mem_11__18_;
   wire Mfifo_psum_M_ffmem_mem_11__19_;
   wire Mfifo_psum_M_ffmem_mem_11__20_;
   wire Mfifo_psum_M_ffmem_mem_11__21_;
   wire Mfifo_psum_M_ffmem_mem_11__22_;
   wire Mfifo_psum_M_ffmem_mem_11__23_;
   wire Mfifo_psum_M_ffmem_mem_11__24_;
   wire Mfifo_psum_M_ffmem_mem_11__25_;
   wire Mfifo_psum_M_ffmem_mem_11__26_;
   wire Mfifo_psum_M_ffmem_mem_11__27_;
   wire Mfifo_psum_M_ffmem_mem_11__28_;
   wire Mfifo_psum_M_ffmem_mem_11__29_;
   wire Mfifo_psum_M_ffmem_mem_11__30_;
   wire Mfifo_psum_M_ffmem_mem_11__31_;
   wire Mfifo_psum_M_ffmem_mem_11__32_;
   wire Mfifo_psum_M_ffmem_mem_11__33_;
   wire Mfifo_psum_M_ffmem_mem_11__34_;
   wire Mfifo_psum_M_ffmem_mem_11__35_;
   wire Mfifo_psum_M_ffmem_mem_11__36_;
   wire Mfifo_psum_M_ffmem_mem_11__37_;
   wire Mfifo_psum_M_ffmem_mem_11__38_;
   wire Mfifo_psum_M_ffmem_mem_11__39_;
   wire Mfifo_psum_M_ffmem_mem_11__40_;
   wire Mfifo_psum_M_ffmem_mem_11__41_;
   wire Mfifo_psum_M_ffmem_mem_10__0_;
   wire Mfifo_psum_M_ffmem_mem_10__1_;
   wire Mfifo_psum_M_ffmem_mem_10__2_;
   wire Mfifo_psum_M_ffmem_mem_10__3_;
   wire Mfifo_psum_M_ffmem_mem_10__4_;
   wire Mfifo_psum_M_ffmem_mem_10__5_;
   wire Mfifo_psum_M_ffmem_mem_10__6_;
   wire Mfifo_psum_M_ffmem_mem_10__7_;
   wire Mfifo_psum_M_ffmem_mem_10__8_;
   wire Mfifo_psum_M_ffmem_mem_10__9_;
   wire Mfifo_psum_M_ffmem_mem_10__10_;
   wire Mfifo_psum_M_ffmem_mem_10__11_;
   wire Mfifo_psum_M_ffmem_mem_10__12_;
   wire Mfifo_psum_M_ffmem_mem_10__13_;
   wire Mfifo_psum_M_ffmem_mem_10__14_;
   wire Mfifo_psum_M_ffmem_mem_10__15_;
   wire Mfifo_psum_M_ffmem_mem_10__16_;
   wire Mfifo_psum_M_ffmem_mem_10__17_;
   wire Mfifo_psum_M_ffmem_mem_10__18_;
   wire Mfifo_psum_M_ffmem_mem_10__19_;
   wire Mfifo_psum_M_ffmem_mem_10__20_;
   wire Mfifo_psum_M_ffmem_mem_10__21_;
   wire Mfifo_psum_M_ffmem_mem_10__22_;
   wire Mfifo_psum_M_ffmem_mem_10__23_;
   wire Mfifo_psum_M_ffmem_mem_10__24_;
   wire Mfifo_psum_M_ffmem_mem_10__25_;
   wire Mfifo_psum_M_ffmem_mem_10__26_;
   wire Mfifo_psum_M_ffmem_mem_10__27_;
   wire Mfifo_psum_M_ffmem_mem_10__28_;
   wire Mfifo_psum_M_ffmem_mem_10__29_;
   wire Mfifo_psum_M_ffmem_mem_10__30_;
   wire Mfifo_psum_M_ffmem_mem_10__31_;
   wire Mfifo_psum_M_ffmem_mem_10__32_;
   wire Mfifo_psum_M_ffmem_mem_10__33_;
   wire Mfifo_psum_M_ffmem_mem_10__34_;
   wire Mfifo_psum_M_ffmem_mem_10__35_;
   wire Mfifo_psum_M_ffmem_mem_10__36_;
   wire Mfifo_psum_M_ffmem_mem_10__37_;
   wire Mfifo_psum_M_ffmem_mem_10__38_;
   wire Mfifo_psum_M_ffmem_mem_10__39_;
   wire Mfifo_psum_M_ffmem_mem_10__40_;
   wire Mfifo_psum_M_ffmem_mem_10__41_;
   wire Mfifo_psum_M_ffmem_mem_9__0_;
   wire Mfifo_psum_M_ffmem_mem_9__1_;
   wire Mfifo_psum_M_ffmem_mem_9__2_;
   wire Mfifo_psum_M_ffmem_mem_9__3_;
   wire Mfifo_psum_M_ffmem_mem_9__4_;
   wire Mfifo_psum_M_ffmem_mem_9__5_;
   wire Mfifo_psum_M_ffmem_mem_9__6_;
   wire Mfifo_psum_M_ffmem_mem_9__7_;
   wire Mfifo_psum_M_ffmem_mem_9__8_;
   wire Mfifo_psum_M_ffmem_mem_9__9_;
   wire Mfifo_psum_M_ffmem_mem_9__10_;
   wire Mfifo_psum_M_ffmem_mem_9__11_;
   wire Mfifo_psum_M_ffmem_mem_9__12_;
   wire Mfifo_psum_M_ffmem_mem_9__13_;
   wire Mfifo_psum_M_ffmem_mem_9__14_;
   wire Mfifo_psum_M_ffmem_mem_9__15_;
   wire Mfifo_psum_M_ffmem_mem_9__16_;
   wire Mfifo_psum_M_ffmem_mem_9__17_;
   wire Mfifo_psum_M_ffmem_mem_9__18_;
   wire Mfifo_psum_M_ffmem_mem_9__19_;
   wire Mfifo_psum_M_ffmem_mem_9__20_;
   wire Mfifo_psum_M_ffmem_mem_9__21_;
   wire Mfifo_psum_M_ffmem_mem_9__22_;
   wire Mfifo_psum_M_ffmem_mem_9__23_;
   wire Mfifo_psum_M_ffmem_mem_9__24_;
   wire Mfifo_psum_M_ffmem_mem_9__25_;
   wire Mfifo_psum_M_ffmem_mem_9__26_;
   wire Mfifo_psum_M_ffmem_mem_9__27_;
   wire Mfifo_psum_M_ffmem_mem_9__28_;
   wire Mfifo_psum_M_ffmem_mem_9__29_;
   wire Mfifo_psum_M_ffmem_mem_9__30_;
   wire Mfifo_psum_M_ffmem_mem_9__31_;
   wire Mfifo_psum_M_ffmem_mem_9__32_;
   wire Mfifo_psum_M_ffmem_mem_9__33_;
   wire Mfifo_psum_M_ffmem_mem_9__34_;
   wire Mfifo_psum_M_ffmem_mem_9__35_;
   wire Mfifo_psum_M_ffmem_mem_9__36_;
   wire Mfifo_psum_M_ffmem_mem_9__37_;
   wire Mfifo_psum_M_ffmem_mem_9__38_;
   wire Mfifo_psum_M_ffmem_mem_9__39_;
   wire Mfifo_psum_M_ffmem_mem_9__40_;
   wire Mfifo_psum_M_ffmem_mem_9__41_;
   wire Mfifo_psum_M_ffmem_mem_8__0_;
   wire Mfifo_psum_M_ffmem_mem_8__1_;
   wire Mfifo_psum_M_ffmem_mem_8__2_;
   wire Mfifo_psum_M_ffmem_mem_8__3_;
   wire Mfifo_psum_M_ffmem_mem_8__4_;
   wire Mfifo_psum_M_ffmem_mem_8__5_;
   wire Mfifo_psum_M_ffmem_mem_8__6_;
   wire Mfifo_psum_M_ffmem_mem_8__7_;
   wire Mfifo_psum_M_ffmem_mem_8__8_;
   wire Mfifo_psum_M_ffmem_mem_8__9_;
   wire Mfifo_psum_M_ffmem_mem_8__10_;
   wire Mfifo_psum_M_ffmem_mem_8__11_;
   wire Mfifo_psum_M_ffmem_mem_8__12_;
   wire Mfifo_psum_M_ffmem_mem_8__13_;
   wire Mfifo_psum_M_ffmem_mem_8__14_;
   wire Mfifo_psum_M_ffmem_mem_8__15_;
   wire Mfifo_psum_M_ffmem_mem_8__16_;
   wire Mfifo_psum_M_ffmem_mem_8__17_;
   wire Mfifo_psum_M_ffmem_mem_8__18_;
   wire Mfifo_psum_M_ffmem_mem_8__19_;
   wire Mfifo_psum_M_ffmem_mem_8__20_;
   wire Mfifo_psum_M_ffmem_mem_8__21_;
   wire Mfifo_psum_M_ffmem_mem_8__22_;
   wire Mfifo_psum_M_ffmem_mem_8__23_;
   wire Mfifo_psum_M_ffmem_mem_8__24_;
   wire Mfifo_psum_M_ffmem_mem_8__25_;
   wire Mfifo_psum_M_ffmem_mem_8__26_;
   wire Mfifo_psum_M_ffmem_mem_8__27_;
   wire Mfifo_psum_M_ffmem_mem_8__28_;
   wire Mfifo_psum_M_ffmem_mem_8__29_;
   wire Mfifo_psum_M_ffmem_mem_8__30_;
   wire Mfifo_psum_M_ffmem_mem_8__31_;
   wire Mfifo_psum_M_ffmem_mem_8__32_;
   wire Mfifo_psum_M_ffmem_mem_8__33_;
   wire Mfifo_psum_M_ffmem_mem_8__34_;
   wire Mfifo_psum_M_ffmem_mem_8__35_;
   wire Mfifo_psum_M_ffmem_mem_8__36_;
   wire Mfifo_psum_M_ffmem_mem_8__37_;
   wire Mfifo_psum_M_ffmem_mem_8__38_;
   wire Mfifo_psum_M_ffmem_mem_8__39_;
   wire Mfifo_psum_M_ffmem_mem_8__40_;
   wire Mfifo_psum_M_ffmem_mem_8__41_;
   wire Mfifo_psum_M_ffmem_mem_7__0_;
   wire Mfifo_psum_M_ffmem_mem_7__1_;
   wire Mfifo_psum_M_ffmem_mem_7__2_;
   wire Mfifo_psum_M_ffmem_mem_7__3_;
   wire Mfifo_psum_M_ffmem_mem_7__4_;
   wire Mfifo_psum_M_ffmem_mem_7__5_;
   wire Mfifo_psum_M_ffmem_mem_7__6_;
   wire Mfifo_psum_M_ffmem_mem_7__7_;
   wire Mfifo_psum_M_ffmem_mem_7__8_;
   wire Mfifo_psum_M_ffmem_mem_7__9_;
   wire Mfifo_psum_M_ffmem_mem_7__10_;
   wire Mfifo_psum_M_ffmem_mem_7__11_;
   wire Mfifo_psum_M_ffmem_mem_7__12_;
   wire Mfifo_psum_M_ffmem_mem_7__13_;
   wire Mfifo_psum_M_ffmem_mem_7__14_;
   wire Mfifo_psum_M_ffmem_mem_7__15_;
   wire Mfifo_psum_M_ffmem_mem_7__16_;
   wire Mfifo_psum_M_ffmem_mem_7__17_;
   wire Mfifo_psum_M_ffmem_mem_7__18_;
   wire Mfifo_psum_M_ffmem_mem_7__19_;
   wire Mfifo_psum_M_ffmem_mem_7__20_;
   wire Mfifo_psum_M_ffmem_mem_7__21_;
   wire Mfifo_psum_M_ffmem_mem_7__22_;
   wire Mfifo_psum_M_ffmem_mem_7__23_;
   wire Mfifo_psum_M_ffmem_mem_7__24_;
   wire Mfifo_psum_M_ffmem_mem_7__25_;
   wire Mfifo_psum_M_ffmem_mem_7__26_;
   wire Mfifo_psum_M_ffmem_mem_7__27_;
   wire Mfifo_psum_M_ffmem_mem_7__28_;
   wire Mfifo_psum_M_ffmem_mem_7__29_;
   wire Mfifo_psum_M_ffmem_mem_7__30_;
   wire Mfifo_psum_M_ffmem_mem_7__31_;
   wire Mfifo_psum_M_ffmem_mem_7__32_;
   wire Mfifo_psum_M_ffmem_mem_7__33_;
   wire Mfifo_psum_M_ffmem_mem_7__34_;
   wire Mfifo_psum_M_ffmem_mem_7__35_;
   wire Mfifo_psum_M_ffmem_mem_7__36_;
   wire Mfifo_psum_M_ffmem_mem_7__37_;
   wire Mfifo_psum_M_ffmem_mem_7__38_;
   wire Mfifo_psum_M_ffmem_mem_7__39_;
   wire Mfifo_psum_M_ffmem_mem_7__40_;
   wire Mfifo_psum_M_ffmem_mem_7__41_;
   wire Mfifo_psum_M_ffmem_mem_6__0_;
   wire Mfifo_psum_M_ffmem_mem_6__1_;
   wire Mfifo_psum_M_ffmem_mem_6__2_;
   wire Mfifo_psum_M_ffmem_mem_6__3_;
   wire Mfifo_psum_M_ffmem_mem_6__4_;
   wire Mfifo_psum_M_ffmem_mem_6__5_;
   wire Mfifo_psum_M_ffmem_mem_6__6_;
   wire Mfifo_psum_M_ffmem_mem_6__7_;
   wire Mfifo_psum_M_ffmem_mem_6__8_;
   wire Mfifo_psum_M_ffmem_mem_6__9_;
   wire Mfifo_psum_M_ffmem_mem_6__10_;
   wire Mfifo_psum_M_ffmem_mem_6__11_;
   wire Mfifo_psum_M_ffmem_mem_6__12_;
   wire Mfifo_psum_M_ffmem_mem_6__13_;
   wire Mfifo_psum_M_ffmem_mem_6__14_;
   wire Mfifo_psum_M_ffmem_mem_6__15_;
   wire Mfifo_psum_M_ffmem_mem_6__16_;
   wire Mfifo_psum_M_ffmem_mem_6__17_;
   wire Mfifo_psum_M_ffmem_mem_6__18_;
   wire Mfifo_psum_M_ffmem_mem_6__19_;
   wire Mfifo_psum_M_ffmem_mem_6__20_;
   wire Mfifo_psum_M_ffmem_mem_6__21_;
   wire Mfifo_psum_M_ffmem_mem_6__22_;
   wire Mfifo_psum_M_ffmem_mem_6__23_;
   wire Mfifo_psum_M_ffmem_mem_6__24_;
   wire Mfifo_psum_M_ffmem_mem_6__25_;
   wire Mfifo_psum_M_ffmem_mem_6__26_;
   wire Mfifo_psum_M_ffmem_mem_6__27_;
   wire Mfifo_psum_M_ffmem_mem_6__28_;
   wire Mfifo_psum_M_ffmem_mem_6__29_;
   wire Mfifo_psum_M_ffmem_mem_6__30_;
   wire Mfifo_psum_M_ffmem_mem_6__31_;
   wire Mfifo_psum_M_ffmem_mem_6__32_;
   wire Mfifo_psum_M_ffmem_mem_6__33_;
   wire Mfifo_psum_M_ffmem_mem_6__34_;
   wire Mfifo_psum_M_ffmem_mem_6__35_;
   wire Mfifo_psum_M_ffmem_mem_6__36_;
   wire Mfifo_psum_M_ffmem_mem_6__37_;
   wire Mfifo_psum_M_ffmem_mem_6__38_;
   wire Mfifo_psum_M_ffmem_mem_6__39_;
   wire Mfifo_psum_M_ffmem_mem_6__40_;
   wire Mfifo_psum_M_ffmem_mem_6__41_;
   wire Mfifo_psum_M_ffmem_mem_5__0_;
   wire Mfifo_psum_M_ffmem_mem_5__1_;
   wire Mfifo_psum_M_ffmem_mem_5__2_;
   wire Mfifo_psum_M_ffmem_mem_5__3_;
   wire Mfifo_psum_M_ffmem_mem_5__4_;
   wire Mfifo_psum_M_ffmem_mem_5__5_;
   wire Mfifo_psum_M_ffmem_mem_5__6_;
   wire Mfifo_psum_M_ffmem_mem_5__7_;
   wire Mfifo_psum_M_ffmem_mem_5__8_;
   wire Mfifo_psum_M_ffmem_mem_5__9_;
   wire Mfifo_psum_M_ffmem_mem_5__10_;
   wire Mfifo_psum_M_ffmem_mem_5__11_;
   wire Mfifo_psum_M_ffmem_mem_5__12_;
   wire Mfifo_psum_M_ffmem_mem_5__13_;
   wire Mfifo_psum_M_ffmem_mem_5__14_;
   wire Mfifo_psum_M_ffmem_mem_5__15_;
   wire Mfifo_psum_M_ffmem_mem_5__16_;
   wire Mfifo_psum_M_ffmem_mem_5__17_;
   wire Mfifo_psum_M_ffmem_mem_5__18_;
   wire Mfifo_psum_M_ffmem_mem_5__19_;
   wire Mfifo_psum_M_ffmem_mem_5__20_;
   wire Mfifo_psum_M_ffmem_mem_5__21_;
   wire Mfifo_psum_M_ffmem_mem_5__22_;
   wire Mfifo_psum_M_ffmem_mem_5__23_;
   wire Mfifo_psum_M_ffmem_mem_5__24_;
   wire Mfifo_psum_M_ffmem_mem_5__25_;
   wire Mfifo_psum_M_ffmem_mem_5__26_;
   wire Mfifo_psum_M_ffmem_mem_5__27_;
   wire Mfifo_psum_M_ffmem_mem_5__28_;
   wire Mfifo_psum_M_ffmem_mem_5__29_;
   wire Mfifo_psum_M_ffmem_mem_5__30_;
   wire Mfifo_psum_M_ffmem_mem_5__31_;
   wire Mfifo_psum_M_ffmem_mem_5__32_;
   wire Mfifo_psum_M_ffmem_mem_5__33_;
   wire Mfifo_psum_M_ffmem_mem_5__34_;
   wire Mfifo_psum_M_ffmem_mem_5__35_;
   wire Mfifo_psum_M_ffmem_mem_5__36_;
   wire Mfifo_psum_M_ffmem_mem_5__37_;
   wire Mfifo_psum_M_ffmem_mem_5__38_;
   wire Mfifo_psum_M_ffmem_mem_5__39_;
   wire Mfifo_psum_M_ffmem_mem_5__40_;
   wire Mfifo_psum_M_ffmem_mem_5__41_;
   wire Mfifo_psum_M_ffmem_mem_4__0_;
   wire Mfifo_psum_M_ffmem_mem_4__1_;
   wire Mfifo_psum_M_ffmem_mem_4__2_;
   wire Mfifo_psum_M_ffmem_mem_4__3_;
   wire Mfifo_psum_M_ffmem_mem_4__4_;
   wire Mfifo_psum_M_ffmem_mem_4__5_;
   wire Mfifo_psum_M_ffmem_mem_4__6_;
   wire Mfifo_psum_M_ffmem_mem_4__7_;
   wire Mfifo_psum_M_ffmem_mem_4__8_;
   wire Mfifo_psum_M_ffmem_mem_4__9_;
   wire Mfifo_psum_M_ffmem_mem_4__10_;
   wire Mfifo_psum_M_ffmem_mem_4__11_;
   wire Mfifo_psum_M_ffmem_mem_4__12_;
   wire Mfifo_psum_M_ffmem_mem_4__13_;
   wire Mfifo_psum_M_ffmem_mem_4__14_;
   wire Mfifo_psum_M_ffmem_mem_4__15_;
   wire Mfifo_psum_M_ffmem_mem_4__16_;
   wire Mfifo_psum_M_ffmem_mem_4__17_;
   wire Mfifo_psum_M_ffmem_mem_4__18_;
   wire Mfifo_psum_M_ffmem_mem_4__19_;
   wire Mfifo_psum_M_ffmem_mem_4__20_;
   wire Mfifo_psum_M_ffmem_mem_4__21_;
   wire Mfifo_psum_M_ffmem_mem_4__22_;
   wire Mfifo_psum_M_ffmem_mem_4__23_;
   wire Mfifo_psum_M_ffmem_mem_4__24_;
   wire Mfifo_psum_M_ffmem_mem_4__25_;
   wire Mfifo_psum_M_ffmem_mem_4__26_;
   wire Mfifo_psum_M_ffmem_mem_4__27_;
   wire Mfifo_psum_M_ffmem_mem_4__28_;
   wire Mfifo_psum_M_ffmem_mem_4__29_;
   wire Mfifo_psum_M_ffmem_mem_4__30_;
   wire Mfifo_psum_M_ffmem_mem_4__31_;
   wire Mfifo_psum_M_ffmem_mem_4__32_;
   wire Mfifo_psum_M_ffmem_mem_4__33_;
   wire Mfifo_psum_M_ffmem_mem_4__34_;
   wire Mfifo_psum_M_ffmem_mem_4__35_;
   wire Mfifo_psum_M_ffmem_mem_4__36_;
   wire Mfifo_psum_M_ffmem_mem_4__37_;
   wire Mfifo_psum_M_ffmem_mem_4__38_;
   wire Mfifo_psum_M_ffmem_mem_4__39_;
   wire Mfifo_psum_M_ffmem_mem_4__40_;
   wire Mfifo_psum_M_ffmem_mem_4__41_;
   wire Mfifo_psum_M_ffmem_mem_3__0_;
   wire Mfifo_psum_M_ffmem_mem_3__1_;
   wire Mfifo_psum_M_ffmem_mem_3__2_;
   wire Mfifo_psum_M_ffmem_mem_3__3_;
   wire Mfifo_psum_M_ffmem_mem_3__4_;
   wire Mfifo_psum_M_ffmem_mem_3__5_;
   wire Mfifo_psum_M_ffmem_mem_3__6_;
   wire Mfifo_psum_M_ffmem_mem_3__7_;
   wire Mfifo_psum_M_ffmem_mem_3__8_;
   wire Mfifo_psum_M_ffmem_mem_3__9_;
   wire Mfifo_psum_M_ffmem_mem_3__10_;
   wire Mfifo_psum_M_ffmem_mem_3__11_;
   wire Mfifo_psum_M_ffmem_mem_3__12_;
   wire Mfifo_psum_M_ffmem_mem_3__13_;
   wire Mfifo_psum_M_ffmem_mem_3__14_;
   wire Mfifo_psum_M_ffmem_mem_3__15_;
   wire Mfifo_psum_M_ffmem_mem_3__16_;
   wire Mfifo_psum_M_ffmem_mem_3__17_;
   wire Mfifo_psum_M_ffmem_mem_3__18_;
   wire Mfifo_psum_M_ffmem_mem_3__19_;
   wire Mfifo_psum_M_ffmem_mem_3__20_;
   wire Mfifo_psum_M_ffmem_mem_3__21_;
   wire Mfifo_psum_M_ffmem_mem_3__22_;
   wire Mfifo_psum_M_ffmem_mem_3__23_;
   wire Mfifo_psum_M_ffmem_mem_3__24_;
   wire Mfifo_psum_M_ffmem_mem_3__25_;
   wire Mfifo_psum_M_ffmem_mem_3__26_;
   wire Mfifo_psum_M_ffmem_mem_3__27_;
   wire Mfifo_psum_M_ffmem_mem_3__28_;
   wire Mfifo_psum_M_ffmem_mem_3__29_;
   wire Mfifo_psum_M_ffmem_mem_3__30_;
   wire Mfifo_psum_M_ffmem_mem_3__31_;
   wire Mfifo_psum_M_ffmem_mem_3__32_;
   wire Mfifo_psum_M_ffmem_mem_3__33_;
   wire Mfifo_psum_M_ffmem_mem_3__34_;
   wire Mfifo_psum_M_ffmem_mem_3__35_;
   wire Mfifo_psum_M_ffmem_mem_3__36_;
   wire Mfifo_psum_M_ffmem_mem_3__37_;
   wire Mfifo_psum_M_ffmem_mem_3__38_;
   wire Mfifo_psum_M_ffmem_mem_3__39_;
   wire Mfifo_psum_M_ffmem_mem_3__40_;
   wire Mfifo_psum_M_ffmem_mem_3__41_;
   wire Mfifo_psum_M_ffmem_mem_2__0_;
   wire Mfifo_psum_M_ffmem_mem_2__1_;
   wire Mfifo_psum_M_ffmem_mem_2__2_;
   wire Mfifo_psum_M_ffmem_mem_2__3_;
   wire Mfifo_psum_M_ffmem_mem_2__4_;
   wire Mfifo_psum_M_ffmem_mem_2__5_;
   wire Mfifo_psum_M_ffmem_mem_2__6_;
   wire Mfifo_psum_M_ffmem_mem_2__7_;
   wire Mfifo_psum_M_ffmem_mem_2__8_;
   wire Mfifo_psum_M_ffmem_mem_2__9_;
   wire Mfifo_psum_M_ffmem_mem_2__10_;
   wire Mfifo_psum_M_ffmem_mem_2__11_;
   wire Mfifo_psum_M_ffmem_mem_2__12_;
   wire Mfifo_psum_M_ffmem_mem_2__13_;
   wire Mfifo_psum_M_ffmem_mem_2__14_;
   wire Mfifo_psum_M_ffmem_mem_2__15_;
   wire Mfifo_psum_M_ffmem_mem_2__16_;
   wire Mfifo_psum_M_ffmem_mem_2__17_;
   wire Mfifo_psum_M_ffmem_mem_2__18_;
   wire Mfifo_psum_M_ffmem_mem_2__19_;
   wire Mfifo_psum_M_ffmem_mem_2__20_;
   wire Mfifo_psum_M_ffmem_mem_2__21_;
   wire Mfifo_psum_M_ffmem_mem_2__22_;
   wire Mfifo_psum_M_ffmem_mem_2__23_;
   wire Mfifo_psum_M_ffmem_mem_2__24_;
   wire Mfifo_psum_M_ffmem_mem_2__25_;
   wire Mfifo_psum_M_ffmem_mem_2__26_;
   wire Mfifo_psum_M_ffmem_mem_2__27_;
   wire Mfifo_psum_M_ffmem_mem_2__28_;
   wire Mfifo_psum_M_ffmem_mem_2__29_;
   wire Mfifo_psum_M_ffmem_mem_2__30_;
   wire Mfifo_psum_M_ffmem_mem_2__31_;
   wire Mfifo_psum_M_ffmem_mem_2__32_;
   wire Mfifo_psum_M_ffmem_mem_2__33_;
   wire Mfifo_psum_M_ffmem_mem_2__34_;
   wire Mfifo_psum_M_ffmem_mem_2__35_;
   wire Mfifo_psum_M_ffmem_mem_2__36_;
   wire Mfifo_psum_M_ffmem_mem_2__37_;
   wire Mfifo_psum_M_ffmem_mem_2__38_;
   wire Mfifo_psum_M_ffmem_mem_2__39_;
   wire Mfifo_psum_M_ffmem_mem_2__40_;
   wire Mfifo_psum_M_ffmem_mem_2__41_;
   wire Mfifo_psum_M_ffmem_mem_1__0_;
   wire Mfifo_psum_M_ffmem_mem_1__1_;
   wire Mfifo_psum_M_ffmem_mem_1__2_;
   wire Mfifo_psum_M_ffmem_mem_1__3_;
   wire Mfifo_psum_M_ffmem_mem_1__4_;
   wire Mfifo_psum_M_ffmem_mem_1__5_;
   wire Mfifo_psum_M_ffmem_mem_1__6_;
   wire Mfifo_psum_M_ffmem_mem_1__7_;
   wire Mfifo_psum_M_ffmem_mem_1__8_;
   wire Mfifo_psum_M_ffmem_mem_1__9_;
   wire Mfifo_psum_M_ffmem_mem_1__10_;
   wire Mfifo_psum_M_ffmem_mem_1__11_;
   wire Mfifo_psum_M_ffmem_mem_1__12_;
   wire Mfifo_psum_M_ffmem_mem_1__13_;
   wire Mfifo_psum_M_ffmem_mem_1__14_;
   wire Mfifo_psum_M_ffmem_mem_1__15_;
   wire Mfifo_psum_M_ffmem_mem_1__16_;
   wire Mfifo_psum_M_ffmem_mem_1__17_;
   wire Mfifo_psum_M_ffmem_mem_1__18_;
   wire Mfifo_psum_M_ffmem_mem_1__19_;
   wire Mfifo_psum_M_ffmem_mem_1__20_;
   wire Mfifo_psum_M_ffmem_mem_1__21_;
   wire Mfifo_psum_M_ffmem_mem_1__22_;
   wire Mfifo_psum_M_ffmem_mem_1__23_;
   wire Mfifo_psum_M_ffmem_mem_1__24_;
   wire Mfifo_psum_M_ffmem_mem_1__25_;
   wire Mfifo_psum_M_ffmem_mem_1__26_;
   wire Mfifo_psum_M_ffmem_mem_1__27_;
   wire Mfifo_psum_M_ffmem_mem_1__28_;
   wire Mfifo_psum_M_ffmem_mem_1__29_;
   wire Mfifo_psum_M_ffmem_mem_1__30_;
   wire Mfifo_psum_M_ffmem_mem_1__31_;
   wire Mfifo_psum_M_ffmem_mem_1__32_;
   wire Mfifo_psum_M_ffmem_mem_1__33_;
   wire Mfifo_psum_M_ffmem_mem_1__34_;
   wire Mfifo_psum_M_ffmem_mem_1__35_;
   wire Mfifo_psum_M_ffmem_mem_1__36_;
   wire Mfifo_psum_M_ffmem_mem_1__37_;
   wire Mfifo_psum_M_ffmem_mem_1__38_;
   wire Mfifo_psum_M_ffmem_mem_1__39_;
   wire Mfifo_psum_M_ffmem_mem_1__40_;
   wire Mfifo_psum_M_ffmem_mem_1__41_;
   wire Mfifo_psum_M_ffmem_mem_0__0_;
   wire Mfifo_psum_M_ffmem_mem_0__1_;
   wire Mfifo_psum_M_ffmem_mem_0__2_;
   wire Mfifo_psum_M_ffmem_mem_0__3_;
   wire Mfifo_psum_M_ffmem_mem_0__4_;
   wire Mfifo_psum_M_ffmem_mem_0__5_;
   wire Mfifo_psum_M_ffmem_mem_0__6_;
   wire Mfifo_psum_M_ffmem_mem_0__7_;
   wire Mfifo_psum_M_ffmem_mem_0__8_;
   wire Mfifo_psum_M_ffmem_mem_0__9_;
   wire Mfifo_psum_M_ffmem_mem_0__10_;
   wire Mfifo_psum_M_ffmem_mem_0__11_;
   wire Mfifo_psum_M_ffmem_mem_0__12_;
   wire Mfifo_psum_M_ffmem_mem_0__13_;
   wire Mfifo_psum_M_ffmem_mem_0__14_;
   wire Mfifo_psum_M_ffmem_mem_0__15_;
   wire Mfifo_psum_M_ffmem_mem_0__16_;
   wire Mfifo_psum_M_ffmem_mem_0__17_;
   wire Mfifo_psum_M_ffmem_mem_0__18_;
   wire Mfifo_psum_M_ffmem_mem_0__19_;
   wire Mfifo_psum_M_ffmem_mem_0__20_;
   wire Mfifo_psum_M_ffmem_mem_0__21_;
   wire Mfifo_psum_M_ffmem_mem_0__22_;
   wire Mfifo_psum_M_ffmem_mem_0__23_;
   wire Mfifo_psum_M_ffmem_mem_0__24_;
   wire Mfifo_psum_M_ffmem_mem_0__25_;
   wire Mfifo_psum_M_ffmem_mem_0__26_;
   wire Mfifo_psum_M_ffmem_mem_0__27_;
   wire Mfifo_psum_M_ffmem_mem_0__28_;
   wire Mfifo_psum_M_ffmem_mem_0__29_;
   wire Mfifo_psum_M_ffmem_mem_0__30_;
   wire Mfifo_psum_M_ffmem_mem_0__31_;
   wire Mfifo_psum_M_ffmem_mem_0__32_;
   wire Mfifo_psum_M_ffmem_mem_0__33_;
   wire Mfifo_psum_M_ffmem_mem_0__34_;
   wire Mfifo_psum_M_ffmem_mem_0__35_;
   wire Mfifo_psum_M_ffmem_mem_0__36_;
   wire Mfifo_psum_M_ffmem_mem_0__37_;
   wire Mfifo_psum_M_ffmem_mem_0__38_;
   wire Mfifo_psum_M_ffmem_mem_0__39_;
   wire Mfifo_psum_M_ffmem_mem_0__40_;
   wire Mfifo_psum_M_ffmem_mem_0__41_;
   wire Mfifo_xin_M_ffmem_mem_15__0_;
   wire Mfifo_xin_M_ffmem_mem_15__1_;
   wire Mfifo_xin_M_ffmem_mem_15__2_;
   wire Mfifo_xin_M_ffmem_mem_15__3_;
   wire Mfifo_xin_M_ffmem_mem_15__4_;
   wire Mfifo_xin_M_ffmem_mem_15__5_;
   wire Mfifo_xin_M_ffmem_mem_15__6_;
   wire Mfifo_xin_M_ffmem_mem_15__7_;
   wire Mfifo_xin_M_ffmem_mem_14__0_;
   wire Mfifo_xin_M_ffmem_mem_14__1_;
   wire Mfifo_xin_M_ffmem_mem_14__2_;
   wire Mfifo_xin_M_ffmem_mem_14__3_;
   wire Mfifo_xin_M_ffmem_mem_14__4_;
   wire Mfifo_xin_M_ffmem_mem_14__5_;
   wire Mfifo_xin_M_ffmem_mem_14__6_;
   wire Mfifo_xin_M_ffmem_mem_14__7_;
   wire Mfifo_xin_M_ffmem_mem_13__0_;
   wire Mfifo_xin_M_ffmem_mem_13__1_;
   wire Mfifo_xin_M_ffmem_mem_13__2_;
   wire Mfifo_xin_M_ffmem_mem_13__3_;
   wire Mfifo_xin_M_ffmem_mem_13__4_;
   wire Mfifo_xin_M_ffmem_mem_13__5_;
   wire Mfifo_xin_M_ffmem_mem_13__6_;
   wire Mfifo_xin_M_ffmem_mem_13__7_;
   wire Mfifo_xin_M_ffmem_mem_12__0_;
   wire Mfifo_xin_M_ffmem_mem_12__1_;
   wire Mfifo_xin_M_ffmem_mem_12__2_;
   wire Mfifo_xin_M_ffmem_mem_12__3_;
   wire Mfifo_xin_M_ffmem_mem_12__4_;
   wire Mfifo_xin_M_ffmem_mem_12__5_;
   wire Mfifo_xin_M_ffmem_mem_12__6_;
   wire Mfifo_xin_M_ffmem_mem_12__7_;
   wire Mfifo_xin_M_ffmem_mem_11__0_;
   wire Mfifo_xin_M_ffmem_mem_11__1_;
   wire Mfifo_xin_M_ffmem_mem_11__2_;
   wire Mfifo_xin_M_ffmem_mem_11__3_;
   wire Mfifo_xin_M_ffmem_mem_11__4_;
   wire Mfifo_xin_M_ffmem_mem_11__5_;
   wire Mfifo_xin_M_ffmem_mem_11__6_;
   wire Mfifo_xin_M_ffmem_mem_11__7_;
   wire Mfifo_xin_M_ffmem_mem_10__0_;
   wire Mfifo_xin_M_ffmem_mem_10__1_;
   wire Mfifo_xin_M_ffmem_mem_10__2_;
   wire Mfifo_xin_M_ffmem_mem_10__3_;
   wire Mfifo_xin_M_ffmem_mem_10__4_;
   wire Mfifo_xin_M_ffmem_mem_10__5_;
   wire Mfifo_xin_M_ffmem_mem_10__6_;
   wire Mfifo_xin_M_ffmem_mem_10__7_;
   wire Mfifo_xin_M_ffmem_mem_9__0_;
   wire Mfifo_xin_M_ffmem_mem_9__1_;
   wire Mfifo_xin_M_ffmem_mem_9__2_;
   wire Mfifo_xin_M_ffmem_mem_9__3_;
   wire Mfifo_xin_M_ffmem_mem_9__4_;
   wire Mfifo_xin_M_ffmem_mem_9__5_;
   wire Mfifo_xin_M_ffmem_mem_9__6_;
   wire Mfifo_xin_M_ffmem_mem_9__7_;
   wire Mfifo_xin_M_ffmem_mem_8__0_;
   wire Mfifo_xin_M_ffmem_mem_8__1_;
   wire Mfifo_xin_M_ffmem_mem_8__2_;
   wire Mfifo_xin_M_ffmem_mem_8__3_;
   wire Mfifo_xin_M_ffmem_mem_8__4_;
   wire Mfifo_xin_M_ffmem_mem_8__5_;
   wire Mfifo_xin_M_ffmem_mem_8__6_;
   wire Mfifo_xin_M_ffmem_mem_8__7_;
   wire Mfifo_xin_M_ffmem_mem_7__0_;
   wire Mfifo_xin_M_ffmem_mem_7__1_;
   wire Mfifo_xin_M_ffmem_mem_7__2_;
   wire Mfifo_xin_M_ffmem_mem_7__3_;
   wire Mfifo_xin_M_ffmem_mem_7__4_;
   wire Mfifo_xin_M_ffmem_mem_7__5_;
   wire Mfifo_xin_M_ffmem_mem_7__6_;
   wire Mfifo_xin_M_ffmem_mem_7__7_;
   wire Mfifo_xin_M_ffmem_mem_6__0_;
   wire Mfifo_xin_M_ffmem_mem_6__1_;
   wire Mfifo_xin_M_ffmem_mem_6__2_;
   wire Mfifo_xin_M_ffmem_mem_6__3_;
   wire Mfifo_xin_M_ffmem_mem_6__4_;
   wire Mfifo_xin_M_ffmem_mem_6__5_;
   wire Mfifo_xin_M_ffmem_mem_6__6_;
   wire Mfifo_xin_M_ffmem_mem_6__7_;
   wire Mfifo_xin_M_ffmem_mem_5__0_;
   wire Mfifo_xin_M_ffmem_mem_5__1_;
   wire Mfifo_xin_M_ffmem_mem_5__2_;
   wire Mfifo_xin_M_ffmem_mem_5__3_;
   wire Mfifo_xin_M_ffmem_mem_5__4_;
   wire Mfifo_xin_M_ffmem_mem_5__5_;
   wire Mfifo_xin_M_ffmem_mem_5__6_;
   wire Mfifo_xin_M_ffmem_mem_5__7_;
   wire Mfifo_xin_M_ffmem_mem_4__0_;
   wire Mfifo_xin_M_ffmem_mem_4__1_;
   wire Mfifo_xin_M_ffmem_mem_4__2_;
   wire Mfifo_xin_M_ffmem_mem_4__3_;
   wire Mfifo_xin_M_ffmem_mem_4__4_;
   wire Mfifo_xin_M_ffmem_mem_4__5_;
   wire Mfifo_xin_M_ffmem_mem_4__6_;
   wire Mfifo_xin_M_ffmem_mem_4__7_;
   wire Mfifo_xin_M_ffmem_mem_3__0_;
   wire Mfifo_xin_M_ffmem_mem_3__1_;
   wire Mfifo_xin_M_ffmem_mem_3__2_;
   wire Mfifo_xin_M_ffmem_mem_3__3_;
   wire Mfifo_xin_M_ffmem_mem_3__4_;
   wire Mfifo_xin_M_ffmem_mem_3__5_;
   wire Mfifo_xin_M_ffmem_mem_3__6_;
   wire Mfifo_xin_M_ffmem_mem_3__7_;
   wire Mfifo_xin_M_ffmem_mem_2__0_;
   wire Mfifo_xin_M_ffmem_mem_2__1_;
   wire Mfifo_xin_M_ffmem_mem_2__2_;
   wire Mfifo_xin_M_ffmem_mem_2__3_;
   wire Mfifo_xin_M_ffmem_mem_2__4_;
   wire Mfifo_xin_M_ffmem_mem_2__5_;
   wire Mfifo_xin_M_ffmem_mem_2__6_;
   wire Mfifo_xin_M_ffmem_mem_2__7_;
   wire Mfifo_xin_M_ffmem_mem_1__0_;
   wire Mfifo_xin_M_ffmem_mem_1__1_;
   wire Mfifo_xin_M_ffmem_mem_1__2_;
   wire Mfifo_xin_M_ffmem_mem_1__3_;
   wire Mfifo_xin_M_ffmem_mem_1__4_;
   wire Mfifo_xin_M_ffmem_mem_1__5_;
   wire Mfifo_xin_M_ffmem_mem_1__6_;
   wire Mfifo_xin_M_ffmem_mem_1__7_;
   wire Mfifo_xin_M_ffmem_mem_0__0_;
   wire Mfifo_xin_M_ffmem_mem_0__1_;
   wire Mfifo_xin_M_ffmem_mem_0__2_;
   wire Mfifo_xin_M_ffmem_mem_0__3_;
   wire Mfifo_xin_M_ffmem_mem_0__4_;
   wire Mfifo_xin_M_ffmem_mem_0__5_;
   wire Mfifo_xin_M_ffmem_mem_0__6_;
   wire Mfifo_xin_M_ffmem_mem_0__7_;
   wire Mfifo_psum_M_rptr_rempty_val;
   wire Mfifo_xin_M_rptr_rempty_val;
   wire Mfifo_xin_M_rptr_N1;
   wire Mfifo_psum_M_wptr_wfull_val;
   wire Mfifo_xin_M_wptr_wfull_val;
   wire Msyncout_synesend_sync2;
   wire Msyncout_synesend_sync1;
   wire Msyncout_synepsum_sync2;
   wire Msyncout_synepsum_sync1;
   wire Msyncout_syneread_sync2;
   wire Msyncout_syneread_sync1;
   wire Msyncin_synsend_sync2;
   wire Msyncin_synsend_sync1;
   wire Msyncin_syncomp_sync2;
   wire Msyncin_syncomp_sync1;
   wire Msyncin_synenable_sync2;
   wire Msyncin_synenable_sync1;
   wire Msyncin_MsynWH_3__synH_sync2;
   wire Msyncin_MsynWH_3__synH_sync1;
   wire Msyncin_MsynWH_3__synW_sync2;
   wire Msyncin_MsynWH_3__synW_sync1;
   wire Msyncin_MsynWH_2__synH_sync2;
   wire Msyncin_MsynWH_2__synH_sync1;
   wire Msyncin_MsynWH_2__synW_sync2;
   wire Msyncin_MsynWH_2__synW_sync1;
   wire Msyncin_MsynWH_1__synH_sync2;
   wire Msyncin_MsynWH_1__synH_sync1;
   wire Msyncin_MsynWH_1__synW_sync2;
   wire Msyncin_MsynWH_1__synW_sync1;
   wire Msyncin_MsynWH_0__synH_sync2;
   wire Msyncin_MsynWH_0__synH_sync1;
   wire Msyncin_MsynWH_0__synW_sync2;
   wire Msyncin_MsynWH_0__synW_sync1;
   wire Msyncin_Msynkxy_1__synky_sync2;
   wire Msyncin_Msynkxy_1__synky_sync1;
   wire Msyncin_Msynkxy_1__synkx_sync2;
   wire Msyncin_Msynkxy_1__synkx_sync1;
   wire Msyncin_Msynkxy_0__synky_sync2;
   wire Msyncin_Msynkxy_0__synky_sync1;
   wire C175_DATA2_0;
   wire C175_DATA2_2;
   wire C175_DATA2_3;
   wire C175_DATA2_4;
   wire C174_DATA2_0;
   wire C174_DATA2_1;
   wire C174_DATA2_2;
   wire C174_DATA2_3;
   wire C174_DATA2_4;
   wire C174_DATA2_5;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1516;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1670;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1749;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1818;
   wire n1819;
   wire n1820;
   wire n1821;
   wire n1822;
   wire n1823;
   wire n1824;
   wire n1825;
   wire n1826;
   wire n1827;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1831;
   wire n1832;
   wire n1833;
   wire n1834;
   wire n1835;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire n2102;
   wire n2103;
   wire n2104;
   wire n2105;
   wire n2106;
   wire n2107;
   wire n2108;
   wire n2109;
   wire n2110;
   wire n2111;
   wire n2112;
   wire n2113;
   wire n2114;
   wire n2115;
   wire n2116;
   wire n2117;
   wire n2118;
   wire n2119;
   wire n2120;
   wire n2121;
   wire n2122;
   wire n2123;
   wire n2124;
   wire n2125;
   wire n2126;
   wire n2127;
   wire n2128;
   wire n2129;
   wire n2130;
   wire n2131;
   wire n2132;
   wire n2133;
   wire n2134;
   wire n2135;
   wire n2136;
   wire n2137;
   wire n2138;
   wire n2139;
   wire n2140;
   wire n2141;
   wire n2142;
   wire n2143;
   wire n2144;
   wire n2145;
   wire n2146;
   wire n2147;
   wire n2148;
   wire n2149;
   wire n2150;
   wire n2151;
   wire n2152;
   wire n2153;
   wire n2154;
   wire n2155;
   wire n2156;
   wire n2157;
   wire n2158;
   wire n2159;
   wire n2160;
   wire n2161;
   wire n2162;
   wire n2163;
   wire n2164;
   wire n2165;
   wire n2166;
   wire n2167;
   wire n2168;
   wire n2169;
   wire n2170;
   wire n2171;
   wire n2172;
   wire n2173;
   wire n2174;
   wire n2175;
   wire n2176;
   wire n2177;
   wire n2178;
   wire n2179;
   wire n2180;
   wire n2181;
   wire n2182;
   wire n2183;
   wire n2184;
   wire n2185;
   wire n2186;
   wire n2187;
   wire n2188;
   wire n2189;
   wire n2190;
   wire n2191;
   wire n2192;
   wire n2193;
   wire n2194;
   wire n2195;
   wire n2196;
   wire n2197;
   wire n2198;
   wire n2199;
   wire n2200;
   wire n2201;
   wire n2202;
   wire n2203;
   wire n2204;
   wire n2205;
   wire n2206;
   wire n2207;
   wire n2208;
   wire n2209;
   wire n2210;
   wire n2211;
   wire n2212;
   wire n2213;
   wire n2214;
   wire n2215;
   wire n2216;
   wire n2217;
   wire n2218;
   wire n2219;
   wire n2220;
   wire n2221;
   wire n2222;
   wire n2223;
   wire n2224;
   wire n2225;
   wire n2226;
   wire n2227;
   wire n2228;
   wire n2229;
   wire n2230;
   wire n2231;
   wire n2232;
   wire n2233;
   wire n2234;
   wire n2235;
   wire n2236;
   wire n2237;
   wire n2238;
   wire n2239;
   wire n2240;
   wire n2241;
   wire n2242;
   wire n2243;
   wire n2244;
   wire n2245;
   wire n2246;
   wire n2247;
   wire n2248;
   wire n2249;
   wire n2250;
   wire n2251;
   wire n2252;
   wire n2253;
   wire n2254;
   wire n2255;
   wire n2256;
   wire n2257;
   wire n2258;
   wire n2259;
   wire n2260;
   wire n2261;
   wire n2262;
   wire n2263;
   wire n2264;
   wire n2265;
   wire n2266;
   wire n2267;
   wire n2268;
   wire n2269;
   wire n2270;
   wire n2271;
   wire n2272;
   wire n2273;
   wire n2274;
   wire n2275;
   wire n2276;
   wire n2277;
   wire n2278;
   wire n2279;
   wire n2280;
   wire n2281;
   wire n2282;
   wire n2283;
   wire n2284;
   wire n2285;
   wire n2286;
   wire n2287;
   wire n2288;
   wire n2289;
   wire n2290;
   wire n2291;
   wire n2292;
   wire n2293;
   wire n2294;
   wire n2295;
   wire n2296;
   wire n2297;
   wire n2298;
   wire n2299;
   wire n2300;
   wire n2301;
   wire n2302;
   wire n2303;
   wire n2304;
   wire n2305;
   wire n2306;
   wire n2307;
   wire n2308;
   wire n2309;
   wire n2310;
   wire n2311;
   wire n2312;
   wire n2313;
   wire n2314;
   wire n2315;
   wire n2316;
   wire n2317;
   wire n2318;
   wire n2319;
   wire n2320;
   wire n2321;
   wire n2322;
   wire n2323;
   wire n2324;
   wire n2325;
   wire n2326;
   wire n2327;
   wire n2328;
   wire n2329;
   wire n2330;
   wire n2331;
   wire n2332;
   wire n2333;
   wire n2334;
   wire n2335;
   wire n2336;
   wire n2337;
   wire n2338;
   wire n2339;
   wire n2340;
   wire n2341;
   wire n2342;
   wire n2343;
   wire n2344;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2361;
   wire n2362;
   wire n2363;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2370;
   wire n2371;
   wire n2372;
   wire n2373;
   wire n2374;
   wire n2375;
   wire n2376;
   wire n2377;
   wire n2378;
   wire n2379;
   wire n2380;
   wire n2381;
   wire n2382;
   wire n2383;
   wire n2384;
   wire n2385;
   wire n2386;
   wire n2387;
   wire n2388;
   wire n2389;
   wire n2390;
   wire n2391;
   wire n2392;
   wire n2393;
   wire n2394;
   wire n2395;
   wire n2396;
   wire n2397;
   wire C2_Z_0;
   wire DP_OP_1205J5_125_5849_n15;
   wire DP_OP_1205J5_125_5849_n14;
   wire DP_OP_1205J5_125_5849_n13;
   wire DP_OP_1205J5_125_5849_n12;
   wire DP_OP_1205J5_125_5849_n7;
   wire DP_OP_1205J5_125_5849_n6;
   wire DP_OP_1205J5_125_5849_n5;
   wire DP_OP_1205J5_125_5849_n4;
   wire DP_OP_1205J5_125_5849_n3;
   wire DP_OP_1205J5_125_5849_n2;
   wire DP_OP_1207J5_130_8771_n12;
   wire DP_OP_1207J5_130_8771_n6;
   wire DP_OP_1207J5_130_8771_n4;
   wire DP_OP_1207J5_130_8771_n3;
   wire DP_OP_1207J5_130_8771_n2;
   wire n2398;
   wire n2399;
   wire n2400;
   wire n2401;
   wire n2402;
   wire n2403;
   wire n2404;
   wire n2405;
   wire n2406;
   wire n2407;
   wire n2408;
   wire n2412;
   wire n2413;
   wire n2414;
   wire n2415;
   wire n2416;
   wire n2417;
   wire n2418;
   wire n2419;
   wire n2420;
   wire n2421;
   wire n2422;
   wire n2423;
   wire n2424;
   wire n2425;
   wire n2426;
   wire n2427;
   wire n2428;
   wire n2429;
   wire n2430;
   wire n2431;
   wire n2432;
   wire n2433;
   wire n2434;
   wire n2435;
   wire n2436;
   wire n2437;
   wire n2438;
   wire n2439;
   wire n2440;
   wire n2441;
   wire n2442;
   wire n2443;
   wire n2444;
   wire n2445;
   wire n2446;
   wire n2447;
   wire n2448;
   wire n2449;
   wire n2450;
   wire n2451;
   wire n2452;
   wire n2453;
   wire n2454;
   wire n2455;
   wire n2456;
   wire n2457;
   wire n2458;
   wire n2459;
   wire n2460;
   wire n2461;
   wire n2462;
   wire n2463;
   wire n2464;
   wire n2465;
   wire n2466;
   wire n2467;
   wire n2468;
   wire n2469;
   wire n2470;
   wire n2471;
   wire n2472;
   wire n2473;
   wire n2474;
   wire n2475;
   wire n2476;
   wire n2477;
   wire n2478;
   wire n2479;
   wire n2480;
   wire n2481;
   wire n2482;
   wire n2483;
   wire n2484;
   wire n2485;
   wire n2486;
   wire n2487;
   wire n2488;
   wire n2489;
   wire n2490;
   wire n2491;
   wire n2492;
   wire n2493;
   wire n2494;
   wire n2495;
   wire n2496;
   wire n2497;
   wire n2498;
   wire n2499;
   wire n2500;
   wire n2501;
   wire n2502;
   wire n2503;
   wire n2504;
   wire n2505;
   wire n2506;
   wire n2507;
   wire n2508;
   wire n2509;
   wire n2510;
   wire n2511;
   wire n2512;
   wire n2513;
   wire n2514;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2525;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2529;
   wire n2530;
   wire n2531;
   wire n2532;
   wire n2533;
   wire n2534;
   wire n2535;
   wire n2536;
   wire n2537;
   wire n2538;
   wire n2539;
   wire n2540;
   wire n2541;
   wire n2542;
   wire n2543;
   wire n2544;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2549;
   wire n2550;
   wire n2551;
   wire n2552;
   wire n2553;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2557;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2561;
   wire n2562;
   wire n2563;
   wire n2564;
   wire n2565;
   wire n2566;
   wire n2567;
   wire n2568;
   wire n2569;
   wire n2570;
   wire n2571;
   wire n2572;
   wire n2573;
   wire n2574;
   wire n2575;
   wire n2576;
   wire n2577;
   wire n2578;
   wire n2579;
   wire n2580;
   wire n2581;
   wire n2582;
   wire n2583;
   wire n2584;
   wire n2585;
   wire n2586;
   wire n2587;
   wire n2588;
   wire n2589;
   wire n2590;
   wire n2591;
   wire n2592;
   wire n2593;
   wire n2594;
   wire n2595;
   wire n2596;
   wire n2597;
   wire n2598;
   wire n2599;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2610;
   wire n2611;
   wire n2612;
   wire n2613;
   wire n2614;
   wire n2615;
   wire n2616;
   wire n2617;
   wire n2618;
   wire n2619;
   wire n2620;
   wire n2621;
   wire n2622;
   wire n2623;
   wire n2624;
   wire n2625;
   wire n2626;
   wire n2627;
   wire n2628;
   wire n2629;
   wire n2630;
   wire n2631;
   wire n2632;
   wire n2633;
   wire n2634;
   wire n2635;
   wire n2636;
   wire n2637;
   wire n2638;
   wire n2639;
   wire n2640;
   wire n2641;
   wire n2642;
   wire n2643;
   wire n2644;
   wire n2645;
   wire n2646;
   wire n2647;
   wire n2648;
   wire n2649;
   wire n2650;
   wire n2651;
   wire n2652;
   wire n2653;
   wire n2654;
   wire n2655;
   wire n2656;
   wire n2657;
   wire n2658;
   wire n2659;
   wire n2660;
   wire n2661;
   wire n2662;
   wire n2663;
   wire n2664;
   wire n2665;
   wire n2666;
   wire n2667;
   wire n2668;
   wire n2669;
   wire n2670;
   wire n2671;
   wire n2672;
   wire n2673;
   wire n2674;
   wire n2675;
   wire n2676;
   wire n2677;
   wire n2678;
   wire n2679;
   wire n2680;
   wire n2681;
   wire n2682;
   wire n2683;
   wire n2684;
   wire n2685;
   wire n2686;
   wire n2687;
   wire n2688;
   wire n2689;
   wire n2690;
   wire n2691;
   wire n2692;
   wire n2693;
   wire n2694;
   wire n2695;
   wire n2696;
   wire n2697;
   wire n2698;
   wire n2699;
   wire n2700;
   wire n2701;
   wire n2702;
   wire n2703;
   wire n2704;
   wire n2705;
   wire n2706;
   wire n2707;
   wire n2708;
   wire n2709;
   wire n2710;
   wire n2711;
   wire n2712;
   wire n2713;
   wire n2714;
   wire n2715;
   wire n2716;
   wire n2717;
   wire n2718;
   wire n2719;
   wire n2720;
   wire n2721;
   wire n2722;
   wire n2723;
   wire n2724;
   wire n2725;
   wire n2726;
   wire n2727;
   wire n2728;
   wire n2729;
   wire n2730;
   wire n2731;
   wire n2732;
   wire n2733;
   wire n2734;
   wire n2735;
   wire n2736;
   wire n2737;
   wire n2738;
   wire n2739;
   wire n2740;
   wire n2741;
   wire n2742;
   wire n2743;
   wire n2744;
   wire n2745;
   wire n2746;
   wire n2747;
   wire n2748;
   wire n2749;
   wire n2750;
   wire n2751;
   wire n2752;
   wire n2753;
   wire n2754;
   wire n2755;
   wire n2756;
   wire n2757;
   wire n2758;
   wire n2759;
   wire n2760;
   wire n2761;
   wire n2762;
   wire n2763;
   wire n2764;
   wire n2765;
   wire n2766;
   wire n2767;
   wire n2768;
   wire n2769;
   wire n2770;
   wire n2771;
   wire n2772;
   wire n2773;
   wire n2774;
   wire n2775;
   wire n2776;
   wire n2777;
   wire n2778;
   wire n2779;
   wire n2780;
   wire n2781;
   wire n2782;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2786;
   wire n2787;
   wire n2788;
   wire n2789;
   wire n2790;
   wire n2791;
   wire n2792;
   wire n2793;
   wire n2794;
   wire n2795;
   wire n2796;
   wire n2797;
   wire n2798;
   wire n2799;
   wire n2800;
   wire n2801;
   wire n2802;
   wire n2803;
   wire n2804;
   wire n2805;
   wire n2806;
   wire n2807;
   wire n2808;
   wire n2809;
   wire n2810;
   wire n2811;
   wire n2812;
   wire n2813;
   wire n2814;
   wire n2815;
   wire n2816;
   wire n2817;
   wire n2818;
   wire n2819;
   wire n2820;
   wire n2821;
   wire n2822;
   wire n2823;
   wire n2824;
   wire n2825;
   wire n2826;
   wire n2827;
   wire n2828;
   wire n2829;
   wire n2830;
   wire n2831;
   wire n2832;
   wire n2833;
   wire n2834;
   wire n2835;
   wire n2836;
   wire n2837;
   wire n2838;
   wire n2839;
   wire n2840;
   wire n2841;
   wire n2842;
   wire n2843;
   wire n2844;
   wire n2845;
   wire n2846;
   wire n2847;
   wire n2848;
   wire n2849;
   wire n2850;
   wire n2851;
   wire n2852;
   wire n2853;
   wire n2854;
   wire n2855;
   wire n2856;
   wire n2857;
   wire n2858;
   wire n2859;
   wire n2860;
   wire n2861;
   wire n2862;
   wire n2863;
   wire n2864;
   wire n2865;
   wire n2866;
   wire n2867;
   wire n2868;
   wire n2869;
   wire n2870;
   wire n2871;
   wire n2872;
   wire n2873;
   wire n2874;
   wire n2875;
   wire n2876;
   wire n2877;
   wire n2878;
   wire n2879;
   wire n2880;
   wire n2881;
   wire n2882;
   wire n2883;
   wire n2884;
   wire n2885;
   wire n2886;
   wire n2887;
   wire n2888;
   wire n2889;
   wire n2890;
   wire n2891;
   wire n2892;
   wire n2893;
   wire n2894;
   wire n2895;
   wire n2896;
   wire n2897;
   wire n2898;
   wire n2899;
   wire n2900;
   wire n2901;
   wire n2902;
   wire n2903;
   wire n2904;
   wire n2905;
   wire n2906;
   wire n2907;
   wire n2908;
   wire n2909;
   wire n2910;
   wire n2911;
   wire n2912;
   wire n2913;
   wire n2914;
   wire n2915;
   wire n2916;
   wire n2917;
   wire n2918;
   wire n2919;
   wire n2920;
   wire n2921;
   wire n2922;
   wire n2923;
   wire n2924;
   wire n2925;
   wire n2926;
   wire n2927;
   wire n2928;
   wire n2929;
   wire n2930;
   wire n2931;
   wire n2932;
   wire n2933;
   wire n2934;
   wire n2935;
   wire n2936;
   wire n2937;
   wire n2938;
   wire n2939;
   wire n2940;
   wire n2941;
   wire n2942;
   wire n2943;
   wire n2944;
   wire n2945;
   wire n2946;
   wire n2947;
   wire n2948;
   wire n2949;
   wire n2950;
   wire n2951;
   wire n2952;
   wire n2953;
   wire n2954;
   wire n2955;
   wire n2956;
   wire n2957;
   wire n2958;
   wire n2959;
   wire n2960;
   wire n2961;
   wire n2962;
   wire n2963;
   wire n2964;
   wire n2965;
   wire n2966;
   wire n2967;
   wire n2968;
   wire n2969;
   wire n2970;
   wire n2971;
   wire n2972;
   wire n2973;
   wire n2974;
   wire n2975;
   wire n2976;
   wire n2977;
   wire n2978;
   wire n2979;
   wire n2980;
   wire n2981;
   wire n2982;
   wire n2983;
   wire n2984;
   wire n2985;
   wire n2986;
   wire n2987;
   wire n2988;
   wire n2989;
   wire n2990;
   wire n2991;
   wire n2992;
   wire n2993;
   wire n2994;
   wire n2995;
   wire n2996;
   wire n2997;
   wire n2998;
   wire n2999;
   wire n3000;
   wire n3001;
   wire n3002;
   wire n3003;
   wire n3004;
   wire n3005;
   wire n3006;
   wire n3007;
   wire n3008;
   wire n3009;
   wire n3010;
   wire n3011;
   wire n3012;
   wire n3013;
   wire n3014;
   wire n3015;
   wire n3016;
   wire n3017;
   wire n3018;
   wire n3019;
   wire n3020;
   wire n3021;
   wire n3022;
   wire n3023;
   wire n3024;
   wire n3025;
   wire n3026;
   wire n3027;
   wire n3028;
   wire n3029;
   wire n3030;
   wire n3031;
   wire n3032;
   wire n3033;
   wire n3034;
   wire n3035;
   wire n3036;
   wire n3037;
   wire n3038;
   wire n3039;
   wire n3040;
   wire n3041;
   wire n3042;
   wire n3043;
   wire n3044;
   wire n3045;
   wire n3046;
   wire n3047;
   wire n3048;
   wire n3049;
   wire n3050;
   wire n3051;
   wire n3052;
   wire n3053;
   wire n3054;
   wire n3055;
   wire n3056;
   wire n3057;
   wire n3058;
   wire n3059;
   wire n3060;
   wire n3061;
   wire n3062;
   wire n3063;
   wire n3064;
   wire n3065;
   wire n3066;
   wire n3067;
   wire n3068;
   wire n3069;
   wire n3070;
   wire n3071;
   wire n3072;
   wire n3073;
   wire n3074;
   wire n3075;
   wire n3076;
   wire n3077;
   wire n3078;
   wire n3079;
   wire n3080;
   wire n3081;
   wire n3082;
   wire n3083;
   wire n3084;
   wire n3085;
   wire n3086;
   wire n3087;
   wire n3088;
   wire n3089;
   wire n3090;
   wire n3091;
   wire n3092;
   wire n3093;
   wire n3094;
   wire n3095;
   wire n3096;
   wire n3097;
   wire n3098;
   wire n3099;
   wire n3100;
   wire n3101;
   wire n3102;
   wire n3103;
   wire n3104;
   wire n3105;
   wire n3106;
   wire n3107;
   wire n3108;
   wire n3109;
   wire n3110;
   wire n3111;
   wire n3112;
   wire n3113;
   wire n3114;
   wire n3115;
   wire n3116;
   wire n3117;
   wire n3118;
   wire n3119;
   wire n3120;
   wire n3121;
   wire n3122;
   wire n3123;
   wire n3124;
   wire n3125;
   wire n3126;
   wire n3127;
   wire n3128;
   wire n3129;
   wire n3130;
   wire n3131;
   wire n3132;
   wire n3133;
   wire n3134;
   wire n3135;
   wire n3136;
   wire n3137;
   wire n3138;
   wire n3139;
   wire n3140;
   wire n3141;
   wire n3142;
   wire n3143;
   wire n3144;
   wire n3145;
   wire n3146;
   wire n3147;
   wire n3148;
   wire n3149;
   wire n3150;
   wire n3151;
   wire n3152;
   wire n3153;
   wire n3154;
   wire n3155;
   wire n3156;
   wire n3157;
   wire n3158;
   wire n3159;
   wire n3160;
   wire n3161;
   wire n3162;
   wire n3163;
   wire n3164;
   wire n3165;
   wire n3166;
   wire n3167;
   wire n3168;
   wire n3169;
   wire n3170;
   wire n3171;
   wire n3172;
   wire n3173;
   wire n3174;
   wire n3175;
   wire n3176;
   wire n3177;
   wire n3178;
   wire n3179;
   wire n3180;
   wire n3181;
   wire n3182;
   wire n3183;
   wire n3184;
   wire n3185;
   wire n3186;
   wire n3187;
   wire n3188;
   wire n3189;
   wire n3190;
   wire n3191;
   wire n3192;
   wire n3193;
   wire n3194;
   wire n3195;
   wire n3196;
   wire n3197;
   wire n3198;
   wire n3199;
   wire n3200;
   wire n3201;
   wire n3202;
   wire n3203;
   wire n3204;
   wire n3205;
   wire n3206;
   wire n3207;
   wire n3208;
   wire n3209;
   wire n3210;
   wire n3211;
   wire n3212;
   wire n3213;
   wire n3214;
   wire n3215;
   wire n3216;
   wire n3217;
   wire n3218;
   wire n3219;
   wire n3220;
   wire n3221;
   wire n3222;
   wire n3223;
   wire n3224;
   wire n3225;
   wire n3226;
   wire n3227;
   wire n3228;
   wire n3229;
   wire n3230;
   wire n3231;
   wire n3232;
   wire n3233;
   wire n3234;
   wire n3235;
   wire n3236;
   wire n3237;
   wire n3238;
   wire n3239;
   wire n3240;
   wire n3241;
   wire n3242;
   wire n3243;
   wire n3244;
   wire n3245;
   wire n3246;
   wire n3247;
   wire n3248;
   wire n3249;
   wire n3250;
   wire n3251;
   wire n3252;
   wire n3253;
   wire n3254;
   wire n3255;
   wire n3256;
   wire n3257;
   wire n3258;
   wire n3259;
   wire n3260;
   wire n3261;
   wire n3262;
   wire n3263;
   wire n3264;
   wire n3265;
   wire n3266;
   wire n3267;
   wire n3268;
   wire n3269;
   wire n3270;
   wire n3271;
   wire n3272;
   wire n3273;
   wire n3274;
   wire n3275;
   wire n3276;
   wire n3277;
   wire n3278;
   wire n3279;
   wire n3280;
   wire n3281;
   wire n3282;
   wire n3283;
   wire n3284;
   wire n3285;
   wire n3286;
   wire n3287;
   wire n3288;
   wire n3289;
   wire n3290;
   wire n3291;
   wire n3292;
   wire n3293;
   wire n3294;
   wire n3295;
   wire n3296;
   wire n3297;
   wire n3298;
   wire n3299;
   wire n3300;
   wire n3301;
   wire n3302;
   wire n3303;
   wire n3304;
   wire n3305;
   wire n3306;
   wire n3307;
   wire n3308;
   wire n3309;
   wire n3310;
   wire n3311;
   wire n3312;
   wire n3313;
   wire n3314;
   wire n3315;
   wire n3316;
   wire n3317;
   wire n3318;
   wire n3319;
   wire n3320;
   wire n3321;
   wire n3322;
   wire n3323;
   wire n3324;
   wire n3325;
   wire n3326;
   wire n3327;
   wire n3328;
   wire n3329;
   wire n3330;
   wire n3331;
   wire n3332;
   wire n3333;
   wire n3334;
   wire n3335;
   wire n3336;
   wire n3337;
   wire n3338;
   wire n3339;
   wire n3340;
   wire n3341;
   wire n3342;
   wire n3343;
   wire n3344;
   wire n3345;
   wire n3346;
   wire n3347;
   wire n3348;
   wire n3349;
   wire n3350;
   wire n3351;
   wire n3352;
   wire n3353;
   wire n3354;
   wire n3355;
   wire n3356;
   wire n3357;
   wire n3358;
   wire n3359;
   wire n3360;
   wire n3361;
   wire n3362;
   wire n3363;
   wire n3364;
   wire n3365;
   wire n3366;
   wire n3367;
   wire n3368;
   wire n3369;
   wire n3370;
   wire n3371;
   wire n3372;
   wire n3373;
   wire n3374;
   wire n3375;
   wire n3376;
   wire n3377;
   wire n3378;
   wire n3379;
   wire n3380;
   wire n3381;
   wire n3382;
   wire n3383;
   wire n3384;
   wire n3385;
   wire n3386;
   wire n3387;
   wire n3388;
   wire n3389;
   wire n3390;
   wire n3391;
   wire n3392;
   wire n3393;
   wire n3394;
   wire n3395;
   wire n3396;
   wire n3397;
   wire n3398;
   wire n3399;
   wire n3400;
   wire n3401;
   wire n3402;
   wire n3403;
   wire n3404;
   wire n3405;
   wire n3406;
   wire n3407;
   wire n3408;
   wire n3409;
   wire n3410;
   wire n3411;
   wire n3412;
   wire n3413;
   wire n3414;
   wire n3415;
   wire n3416;
   wire n3417;
   wire n3418;
   wire n3419;
   wire n3420;
   wire n3421;
   wire n3422;
   wire n3423;
   wire n3424;
   wire n3425;
   wire n3426;
   wire n3427;
   wire n3428;
   wire n3429;
   wire n3430;
   wire n3431;
   wire n3432;
   wire n3433;
   wire n3434;
   wire n3435;
   wire n3436;
   wire n3437;
   wire n3438;
   wire n3439;
   wire n3440;
   wire n3441;
   wire n3442;
   wire n3443;
   wire n3444;
   wire n3445;
   wire n3446;
   wire n3447;
   wire n3448;
   wire n3449;
   wire n3450;
   wire n3451;
   wire n3452;
   wire n3453;
   wire n3454;
   wire n3455;
   wire n3456;
   wire n3457;
   wire n3458;
   wire n3459;
   wire n3460;
   wire n3461;
   wire n3462;
   wire n3463;
   wire n3464;
   wire n3465;
   wire n3466;
   wire n3467;
   wire n3468;
   wire n3469;
   wire n3470;
   wire n3471;
   wire n3472;
   wire n3473;
   wire n3474;
   wire n3475;
   wire n3476;
   wire n3477;
   wire n3478;
   wire n3479;
   wire n3480;
   wire n3481;
   wire n3482;
   wire n3483;
   wire n3484;
   wire n3485;
   wire n3486;
   wire n3487;
   wire n3488;
   wire n3489;
   wire n3490;
   wire n3491;
   wire n3492;
   wire n3493;
   wire n3494;
   wire n3495;
   wire n3496;
   wire n3497;
   wire n3498;
   wire n3499;
   wire n3500;
   wire n3501;
   wire n3502;
   wire n3503;
   wire n3504;
   wire n3505;
   wire n3506;
   wire n3507;
   wire n3508;
   wire n3509;
   wire n3510;
   wire n3511;
   wire n3512;
   wire n3513;
   wire n3514;
   wire n3515;
   wire n3516;
   wire n3517;
   wire n3518;
   wire n3519;
   wire n3520;
   wire n3521;
   wire n3522;
   wire n3523;
   wire n3524;
   wire n3525;
   wire n3526;
   wire n3527;
   wire n3528;
   wire n3529;
   wire n3530;
   wire n3531;
   wire n3532;
   wire n3533;
   wire n3534;
   wire n3535;
   wire n3536;
   wire n3537;
   wire n3538;
   wire n3539;
   wire n3540;
   wire n3541;
   wire n3542;
   wire n3543;
   wire n3544;
   wire n3545;
   wire n3546;
   wire n3547;
   wire n3548;
   wire n3549;
   wire n3550;
   wire n3551;
   wire n3552;
   wire n3553;
   wire n3554;
   wire n3555;
   wire n3556;
   wire n3557;
   wire n3558;
   wire n3559;
   wire n3560;
   wire n3561;
   wire n3562;
   wire n3563;
   wire n3564;
   wire n3565;
   wire n3566;
   wire n3567;
   wire n3568;
   wire n3569;
   wire n3570;
   wire n3571;
   wire n3572;
   wire n3573;
   wire n3574;
   wire n3575;
   wire n3576;
   wire n3577;
   wire n3578;
   wire n3579;
   wire n3580;
   wire n3581;
   wire n3582;
   wire n3583;
   wire n3584;
   wire n3585;
   wire n3586;
   wire n3587;
   wire n3588;
   wire n3589;
   wire n3590;
   wire n3591;
   wire n3592;
   wire n3593;
   wire n3594;
   wire n3595;
   wire n3596;
   wire n3597;
   wire n3598;
   wire n3599;
   wire n3600;
   wire n3601;
   wire n3602;
   wire n3603;
   wire n3604;
   wire n3605;
   wire n3606;
   wire n3607;
   wire n3608;
   wire n3609;
   wire n3610;
   wire n3611;
   wire n3612;
   wire n3613;
   wire n3614;
   wire n3615;
   wire n3616;
   wire n3617;
   wire n3618;
   wire n3619;
   wire n3620;
   wire n3621;
   wire n3622;
   wire n3623;
   wire n3624;
   wire n3625;
   wire n3626;
   wire n3627;
   wire n3628;
   wire n3629;
   wire n3630;
   wire n3631;
   wire n3632;
   wire n3633;
   wire n3634;
   wire n3635;
   wire n3636;
   wire n3637;
   wire n3638;
   wire n3639;
   wire n3640;
   wire n3641;
   wire n3642;
   wire n3643;
   wire n3644;
   wire n3645;
   wire n3646;
   wire n3647;
   wire n3648;
   wire n3649;
   wire n3650;
   wire n3651;
   wire n3652;
   wire n3653;
   wire n3654;
   wire n3655;
   wire n3656;
   wire n3657;
   wire n3658;
   wire n3659;
   wire n3660;
   wire n3661;
   wire n3662;
   wire n3663;
   wire n3664;
   wire n3665;
   wire n3666;
   wire n3667;
   wire n3668;
   wire n3669;
   wire n3670;
   wire n3671;
   wire n3672;
   wire n3673;
   wire n3674;
   wire n3675;
   wire n3676;
   wire n3677;
   wire n3678;
   wire n3679;
   wire n3680;
   wire n3681;
   wire n3682;
   wire n3683;
   wire n3684;
   wire n3685;
   wire n3686;
   wire n3687;
   wire n3688;
   wire n3689;
   wire n3690;
   wire n3691;
   wire n3692;
   wire n3693;
   wire n3694;
   wire n3695;
   wire n3696;
   wire n3697;
   wire n3698;
   wire n3699;
   wire n3700;
   wire n3701;
   wire n3702;
   wire n3703;
   wire n3704;
   wire n3705;
   wire n3706;
   wire n3707;
   wire n3708;
   wire n3709;
   wire n3710;
   wire n3711;
   wire n3712;
   wire n3713;
   wire n3714;
   wire n3715;
   wire n3716;
   wire n3717;
   wire n3718;
   wire n3719;
   wire n3720;
   wire n3721;
   wire n3722;
   wire n3723;
   wire n3724;
   wire n3725;
   wire n3726;
   wire n3727;
   wire n3728;
   wire n3729;
   wire n3730;
   wire n3731;
   wire n3732;
   wire n3733;
   wire n3734;
   wire n3735;
   wire n3736;
   wire n3737;
   wire n3738;
   wire n3739;
   wire n3740;
   wire n3741;
   wire n3742;
   wire n3743;
   wire n3744;
   wire n3745;
   wire n3746;
   wire n3747;
   wire n3748;
   wire n3749;
   wire n3750;
   wire n3751;
   wire n3752;
   wire n3753;
   wire n3754;
   wire n3755;
   wire n3756;
   wire n3757;
   wire n3758;
   wire n3759;
   wire n3760;
   wire n3761;
   wire n3762;
   wire n3763;
   wire n3764;
   wire n3765;
   wire n3766;
   wire n3767;
   wire n3768;
   wire n3769;
   wire n3770;
   wire n3771;
   wire n3772;
   wire n3773;
   wire n3774;
   wire n3775;
   wire n3776;
   wire n3777;
   wire n3778;
   wire n3779;
   wire n3780;
   wire n3781;
   wire n3782;
   wire n3783;
   wire n3784;
   wire n3785;
   wire n3786;
   wire n3787;
   wire n3788;
   wire n3789;
   wire n3790;
   wire n3791;
   wire n3792;
   wire n3793;
   wire n3794;
   wire n3795;
   wire n3796;
   wire n3797;
   wire n3798;
   wire n3799;
   wire n3800;
   wire n3801;
   wire n3802;
   wire n3803;
   wire n3805;
   wire n3806;
   wire n3807;
   wire n3808;
   wire n3809;
   wire n3810;
   wire n3811;
   wire n3812;
   wire n3813;
   wire n3814;
   wire n3815;
   wire n3816;
   wire n3817;
   wire n3818;
   wire n3819;
   wire n3820;
   wire n3821;
   wire n3822;
   wire n3823;
   wire n3824;
   wire n3825;
   wire n3826;
   wire n3827;
   wire n3828;
   wire n3829;
   wire n3830;
   wire n3831;
   wire n3832;
   wire n3833;
   wire n3834;
   wire n3835;
   wire n3836;
   wire n3837;
   wire n3838;
   wire n3839;
   wire n3840;
   wire n3841;
   wire n3842;
   wire n3843;
   wire [1:0] c_kx;
   wire [1:0] c_ky;
   wire [1:0] c_k_cin;
   wire [3:0] c_cout;
   wire [6:0] x_addr;
   wire [3:0] wen_x_reg;
   wire [2:0] count_k;
   wire [5:0] psum_addr;
   wire [1:0] sel_reg;
   wire [1:0] int_kx;
   wire [1:0] int_ky;
   wire [3:0] int_W;
   wire [3:0] int_H;
   wire [7:0] int_coe;
   wire [7:0] int_xin;
   wire [127:0] coe_out;
   wire [7:0] xin1;
   wire [7:0] xin2;
   wire [7:0] xin3;
   wire [7:0] xin4;
   wire [303:0] psum_o1;
   wire [303:0] psum_o2;
   wire [303:0] psum_o3;
   wire [303:0] psum_o4;
   wire [20:0] psum1_o1;
   wire [20:0] psum1_o2;
   wire [20:0] psum1_o3;
   wire [20:0] psum1_o4;
   wire [20:0] psum2_o1;
   wire [20:0] psum2_o2;
   wire [20:0] psum2_o3;
   wire [20:0] psum2_o4;
   wire [20:0] psum3_o1;
   wire [20:0] psum3_o2;
   wire [20:0] psum3_o3;
   wire [20:0] psum3_o4;
   wire [20:0] psum4_o1;
   wire [20:0] psum4_o2;
   wire [20:0] psum4_o3;
   wire [20:0] psum4_o4;
   wire [20:0] psum1_reg1;
   wire [20:0] psum1_reg2;
   wire [20:0] psum1_reg3;
   wire [20:0] psum1_reg4;
   wire [20:0] psum2_reg1;
   wire [20:0] psum2_reg2;
   wire [20:0] psum2_reg3;
   wire [20:0] psum2_reg4;
   wire [20:0] psum3_reg1;
   wire [20:0] psum3_reg2;
   wire [20:0] psum3_reg3;
   wire [20:0] psum3_reg4;
   wire [20:0] psum4_reg1;
   wire [20:0] psum4_reg2;
   wire [20:0] psum4_reg3;
   wire [20:0] psum4_reg4;
   wire [4:0] Mfifo_coe_wq2_rptr;
   wire [4:0] Mfifo_coe_wptr;
   wire [4:0] Mfifo_coe_rq2_wptr;
   wire [4:0] Mfifo_coe_rptr;
   wire [3:0] Mfifo_coe_raddr;
   wire [3:0] Mfifo_coe_waddr;
   wire [4:0] Mfifo_psum_wq2_rptr;
   wire [4:0] Mfifo_psum_wptr;
   wire [4:0] Mfifo_psum_rq2_wptr;
   wire [4:0] Mfifo_psum_rptr;
   wire [3:0] Mfifo_psum_raddr;
   wire [3:0] Mfifo_psum_waddr;
   wire [4:0] Mfifo_xin_wq2_rptr;
   wire [4:0] Mfifo_xin_wptr;
   wire [4:0] Mfifo_xin_rq2_wptr;
   wire [4:0] Mfifo_xin_rptr;
   wire [3:0] Mfifo_xin_raddr;
   wire [3:0] Mfifo_xin_waddr;
   wire [2:0] Mcntl_Mcntl_current_state;
   wire [3:2] Mcntl_Mcntldata_c_p_W;
   wire [1:0] Mcntl_Mcntldata_c_p_cin;
   wire [3:0] Mcntl_Mcntldata_c_p_H;
   wire [1:0] Mcntl_Mcntldata_c_p_wd4;
   wire [2:1] Mcntl_Mcntldata_c_p_cout;
   wire [1:0] Mcntl_Mcntldata_count;
   wire [1:0] Mcntl_Mcntldata_c_W_r4;
   wire [3:0] Mcntl_Mcntldata_c_x_H;
   wire [1:0] Mcntl_Mcntldata_c_W_d4;
   wire [1:0] Mcntl_Mcntldata_c_x_cin;
   wire [1:0] Mcntl_Mcntldata_c_cin;
   wire [3:0] Mcntl_Mcntldata_x_H_reg;
   wire [3:0] Mcntl_Mcntldata_x_W_reg;
   wire [1:0] Mcntl_Mcntldata_ky_reg;
   wire [1:0] Mcntl_Mcntldata_kx_reg;
   wire [3:0] Mfifo_coe_M_rptr_rgraynext;
   wire [4:0] Mfifo_coe_M_rptr_rbinnext;
   wire [3:0] Mfifo_coe_M_wptr_wgraynext;
   wire [4:0] Mfifo_coe_M_wptr_wbinnext;
   wire [4:0] Mfifo_coe_M_r2w_wq3;
   wire [4:0] Mfifo_coe_M_r2w_wq2;
   wire [4:0] Mfifo_coe_M_w2r_rq3;
   wire [4:0] Mfifo_coe_M_w2r_rq2;
   wire [3:0] Mfifo_psum_M_rptr_rgraynext;
   wire [4:0] Mfifo_psum_M_rptr_rbinnext;
   wire [3:0] Mfifo_xin_M_rptr_rgraynext;
   wire [4:0] Mfifo_xin_M_rptr_rbinnext;
   wire [3:0] Mfifo_psum_M_wptr_wgraynext;
   wire [4:0] Mfifo_psum_M_wptr_wbinnext;
   wire [3:0] Mfifo_xin_M_wptr_wgraynext;
   wire [4:0] Mfifo_xin_M_wptr_wbinnext;
   wire [4:0] Mfifo_psum_M_r2w_wq3;
   wire [4:0] Mfifo_psum_M_r2w_wq2;
   wire [4:0] Mfifo_xin_M_r2w_wq3;
   wire [4:0] Mfifo_xin_M_r2w_wq2;
   wire [4:0] Mfifo_psum_M_w2r_rq3;
   wire [4:0] Mfifo_psum_M_w2r_rq2;
   wire [4:0] Mfifo_xin_M_w2r_rq3;
   wire [4:0] Mfifo_xin_M_w2r_rq2;

   // Module instantiations
   Reg_coe_ary_mini MRegm (
	.coe_out(coe_out),
	.coe_in(int_coe),
	.kx(c_kx),
	.ky(c_ky),
	.cin(c_k_cin),
	.cout(c_cout),
	.write(wen_coe),
	.clk(int_clk),
	.rst_n(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_x_block MRegx (
	.xin1(xin1),
	.xin2(xin2),
	.xin3(xin3),
	.xin4(xin4),
	.int_xin(int_xin),
	.wen_x_reg(wen_x_reg),
	.wen_x(wen_x),
	.x_addr(x_addr),
	.int_clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Pre_mux_ary_b MPre_mux_a (
	.psum_o1(psum_o1),
	.psum_o2(psum_o2),
	.psum_o3(psum_o3),
	.psum_o4(psum_o4),
	.xin1(xin1),
	.xin2(xin2),
	.xin3(xin3),
	.xin4(xin4),
	.coein(coe_out),
	.adden(adden),
	.xen1(xen1),
	.xen4(xen4),
	.sel_xen4({ n2397,
		n2396 }),
	.clk(int_clk),
	.rst_n(int_rst_n),
	.coen(coen), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   PsumAdd_block MPsumadd (
	.psum_o1(psum_o1),
	.psum_o2(psum_o2),
	.psum_o3(psum_o3),
	.psum_o4(psum_o4),
	.psum1_o1(psum1_o1),
	.psum1_o2(psum1_o2),
	.psum1_o3(psum1_o3),
	.psum1_o4(psum1_o4),
	.psum2_o1(psum2_o1),
	.psum2_o2(psum2_o2),
	.psum2_o3(psum2_o3),
	.psum2_o4(psum2_o4),
	.psum3_o1(psum3_o1),
	.psum3_o2(psum3_o2),
	.psum3_o3(psum3_o3),
	.psum3_o4(psum3_o4),
	.psum4_o1(psum4_o1),
	.psum4_o2(psum4_o2),
	.psum4_o3(psum4_o3),
	.psum4_o4(psum4_o4),
	.psum1_reg1(psum1_reg1),
	.psum1_reg2(psum1_reg2),
	.psum1_reg3(psum1_reg3),
	.psum1_reg4(psum1_reg4),
	.psum2_reg1(psum2_reg1),
	.psum2_reg2(psum2_reg2),
	.psum2_reg3(psum2_reg3),
	.psum2_reg4(psum2_reg4),
	.psum3_reg1(psum3_reg1),
	.psum3_reg2(psum3_reg2),
	.psum3_reg3(psum3_reg3),
	.psum3_reg4(psum3_reg4),
	.psum4_reg1(psum4_reg1),
	.psum4_reg2(psum4_reg2),
	.psum4_reg3(psum4_reg3),
	.psum4_reg4(psum4_reg4),
	.count_k({ count_k[2],
		count_k[1],
		1'b0 }),
	.adden_sec(adden_sec),
	.int_clk(int_clk),
	.int_rst_n(int_rst_n),
	.kernel_end_BAR(n3839), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_0__synkx_sync2_reg (
	.Q(Msyncin_Msynkxy_0__synkx_sync2),
	.CK(int_clk),
	.D(ext_kx[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_0__synkx_sync1_reg (
	.Q(Msyncin_Msynkxy_0__synkx_sync1),
	.CK(int_clk),
	.D(Msyncin_Msynkxy_0__synkx_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_0__synkx_synced_reg (
	.Q(int_kx[0]),
	.CK(int_clk),
	.D(Msyncin_Msynkxy_0__synkx_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_rptr_rptr_reg_0_ (
	.Q(Mfifo_coe_rptr[0]),
	.CK(int_clk),
	.D(Mfifo_coe_M_rptr_rgraynext[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_rptr_rptr_reg_1_ (
	.Q(Mfifo_coe_rptr[1]),
	.CK(int_clk),
	.D(Mfifo_coe_M_rptr_rgraynext[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_rptr_rptr_reg_2_ (
	.Q(Mfifo_coe_rptr[2]),
	.CK(int_clk),
	.D(Mfifo_coe_M_rptr_rgraynext[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_rptr_rptr_reg_3_ (
	.Q(Mfifo_coe_rptr[3]),
	.CK(int_clk),
	.D(Mfifo_coe_M_rptr_rgraynext[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_rptr_rptr_reg_4_ (
	.Q(Mfifo_coe_rptr[4]),
	.CK(int_clk),
	.D(Mfifo_coe_M_rptr_rbinnext[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_rptr_rbin_reg_0_ (
	.Q(Mfifo_coe_raddr[0]),
	.CK(int_clk),
	.D(Mfifo_coe_M_rptr_rbinnext[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_rptr_rbin_reg_1_ (
	.Q(Mfifo_coe_raddr[1]),
	.CK(int_clk),
	.D(Mfifo_coe_M_rptr_rbinnext[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_rptr_rbin_reg_2_ (
	.Q(Mfifo_coe_raddr[2]),
	.CK(int_clk),
	.D(Mfifo_coe_M_rptr_rbinnext[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_rptr_rbin_reg_3_ (
	.Q(Mfifo_coe_raddr[3]),
	.CK(int_clk),
	.D(Mfifo_coe_M_rptr_rbinnext[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_wptr_wptr_reg_0_ (
	.Q(Mfifo_coe_wptr[0]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_wptr_wgraynext[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_wptr_wptr_reg_1_ (
	.Q(Mfifo_coe_wptr[1]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_wptr_wgraynext[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_wptr_wptr_reg_2_ (
	.Q(Mfifo_coe_wptr[2]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_wptr_wgraynext[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_wptr_wptr_reg_3_ (
	.Q(Mfifo_coe_wptr[3]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_wptr_wgraynext[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_wptr_wptr_reg_4_ (
	.Q(Mfifo_coe_wptr[4]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_wptr_wbinnext[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_wptr_wbin_reg_0_ (
	.Q(Mfifo_coe_waddr[0]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_wptr_wbinnext[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_wptr_wbin_reg_1_ (
	.Q(Mfifo_coe_waddr[1]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_wptr_wbinnext[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_wptr_wbin_reg_2_ (
	.Q(Mfifo_coe_waddr[2]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_wptr_wbinnext[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_wptr_wbin_reg_3_ (
	.Q(Mfifo_coe_waddr[3]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_wptr_wbinnext[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq3_reg_0_ (
	.Q(Mfifo_coe_M_r2w_wq3[0]),
	.CK(ext_clk),
	.D(Mfifo_coe_rptr[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq2_reg_0_ (
	.Q(Mfifo_coe_M_r2w_wq2[0]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_r2w_wq3[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq2_rptr_reg_0_ (
	.Q(Mfifo_coe_wq2_rptr[0]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_r2w_wq2[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq3_reg_1_ (
	.Q(Mfifo_coe_M_r2w_wq3[1]),
	.CK(ext_clk),
	.D(Mfifo_coe_rptr[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq2_reg_1_ (
	.Q(Mfifo_coe_M_r2w_wq2[1]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_r2w_wq3[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq2_rptr_reg_1_ (
	.Q(Mfifo_coe_wq2_rptr[1]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_r2w_wq2[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq3_reg_2_ (
	.Q(Mfifo_coe_M_r2w_wq3[2]),
	.CK(ext_clk),
	.D(Mfifo_coe_rptr[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq2_reg_2_ (
	.Q(Mfifo_coe_M_r2w_wq2[2]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_r2w_wq3[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq2_rptr_reg_2_ (
	.Q(Mfifo_coe_wq2_rptr[2]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_r2w_wq2[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq3_reg_3_ (
	.Q(Mfifo_coe_M_r2w_wq3[3]),
	.CK(ext_clk),
	.D(Mfifo_coe_rptr[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq2_reg_3_ (
	.Q(Mfifo_coe_M_r2w_wq2[3]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_r2w_wq3[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq2_rptr_reg_3_ (
	.Q(Mfifo_coe_wq2_rptr[3]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_r2w_wq2[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq3_reg_4_ (
	.Q(Mfifo_coe_M_r2w_wq3[4]),
	.CK(ext_clk),
	.D(Mfifo_coe_rptr[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq2_reg_4_ (
	.Q(Mfifo_coe_M_r2w_wq2[4]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_r2w_wq3[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_r2w_wq2_rptr_reg_4_ (
	.Q(Mfifo_coe_wq2_rptr[4]),
	.CK(ext_clk),
	.D(Mfifo_coe_M_r2w_wq2[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_wptr_wfull_reg (
	.Q(n3845),
	.CK(ext_clk),
	.D(Mfifo_coe_M_wptr_wfull_val),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq3_reg_0_ (
	.Q(Mfifo_coe_M_w2r_rq3[0]),
	.CK(int_clk),
	.D(Mfifo_coe_wptr[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq2_reg_0_ (
	.Q(Mfifo_coe_M_w2r_rq2[0]),
	.CK(int_clk),
	.D(Mfifo_coe_M_w2r_rq3[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq2_wptr_reg_0_ (
	.Q(Mfifo_coe_rq2_wptr[0]),
	.CK(int_clk),
	.D(Mfifo_coe_M_w2r_rq2[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq3_reg_1_ (
	.Q(Mfifo_coe_M_w2r_rq3[1]),
	.CK(int_clk),
	.D(Mfifo_coe_wptr[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq2_reg_1_ (
	.Q(Mfifo_coe_M_w2r_rq2[1]),
	.CK(int_clk),
	.D(Mfifo_coe_M_w2r_rq3[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq2_wptr_reg_1_ (
	.Q(Mfifo_coe_rq2_wptr[1]),
	.CK(int_clk),
	.D(Mfifo_coe_M_w2r_rq2[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq3_reg_2_ (
	.Q(Mfifo_coe_M_w2r_rq3[2]),
	.CK(int_clk),
	.D(Mfifo_coe_wptr[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq2_reg_2_ (
	.Q(Mfifo_coe_M_w2r_rq2[2]),
	.CK(int_clk),
	.D(Mfifo_coe_M_w2r_rq3[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq2_wptr_reg_2_ (
	.Q(Mfifo_coe_rq2_wptr[2]),
	.CK(int_clk),
	.D(Mfifo_coe_M_w2r_rq2[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq3_reg_3_ (
	.Q(Mfifo_coe_M_w2r_rq3[3]),
	.CK(int_clk),
	.D(Mfifo_coe_wptr[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq2_reg_3_ (
	.Q(Mfifo_coe_M_w2r_rq2[3]),
	.CK(int_clk),
	.D(Mfifo_coe_M_w2r_rq3[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq2_wptr_reg_3_ (
	.Q(Mfifo_coe_rq2_wptr[3]),
	.CK(int_clk),
	.D(Mfifo_coe_M_w2r_rq2[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq3_reg_4_ (
	.Q(Mfifo_coe_M_w2r_rq3[4]),
	.CK(int_clk),
	.D(Mfifo_coe_wptr[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq2_reg_4_ (
	.Q(Mfifo_coe_M_w2r_rq2[4]),
	.CK(int_clk),
	.D(Mfifo_coe_M_w2r_rq3[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_coe_M_w2r_rq2_wptr_reg_4_ (
	.Q(Mfifo_coe_rq2_wptr[4]),
	.CK(int_clk),
	.D(Mfifo_coe_M_w2r_rq2[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_rptr_rptr_reg_0_ (
	.Q(Mfifo_psum_rptr[0]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_rptr_rgraynext[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_rptr_rptr_reg_1_ (
	.Q(Mfifo_psum_rptr[1]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_rptr_rgraynext[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_rptr_rptr_reg_2_ (
	.Q(Mfifo_psum_rptr[2]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_rptr_rgraynext[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_rptr_rptr_reg_3_ (
	.Q(Mfifo_psum_rptr[3]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_rptr_rgraynext[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_rptr_rptr_reg_4_ (
	.Q(Mfifo_psum_rptr[4]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_rptr_rbinnext[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_rptr_rbin_reg_0_ (
	.Q(Mfifo_psum_raddr[0]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_rptr_rbinnext[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_rptr_rbin_reg_1_ (
	.Q(Mfifo_psum_raddr[1]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_rptr_rbinnext[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_rptr_rbin_reg_2_ (
	.Q(Mfifo_psum_raddr[2]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_rptr_rbinnext[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_rptr_rptr_reg_0_ (
	.Q(Mfifo_xin_rptr[0]),
	.CK(int_clk),
	.D(Mfifo_xin_M_rptr_rgraynext[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_rptr_rptr_reg_1_ (
	.Q(Mfifo_xin_rptr[1]),
	.CK(int_clk),
	.D(Mfifo_xin_M_rptr_rgraynext[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_rptr_rptr_reg_2_ (
	.Q(Mfifo_xin_rptr[2]),
	.CK(int_clk),
	.D(Mfifo_xin_M_rptr_rgraynext[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_rptr_rptr_reg_3_ (
	.Q(Mfifo_xin_rptr[3]),
	.CK(int_clk),
	.D(Mfifo_xin_M_rptr_rgraynext[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_rptr_rptr_reg_4_ (
	.Q(Mfifo_xin_rptr[4]),
	.CK(int_clk),
	.D(Mfifo_xin_M_rptr_rbinnext[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_rptr_rbin_reg_0_ (
	.Q(Mfifo_xin_raddr[0]),
	.CK(int_clk),
	.D(Mfifo_xin_M_rptr_rbinnext[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_rptr_rbin_reg_1_ (
	.Q(Mfifo_xin_raddr[1]),
	.CK(int_clk),
	.D(Mfifo_xin_M_rptr_rbinnext[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_rptr_rbin_reg_3_ (
	.Q(Mfifo_xin_raddr[3]),
	.CK(int_clk),
	.D(Mfifo_xin_M_rptr_rbinnext[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_wptr_wptr_reg_0_ (
	.Q(Mfifo_psum_wptr[0]),
	.CK(int_clk),
	.D(Mfifo_psum_M_wptr_wgraynext[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_wptr_wptr_reg_1_ (
	.Q(Mfifo_psum_wptr[1]),
	.CK(int_clk),
	.D(Mfifo_psum_M_wptr_wgraynext[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_wptr_wptr_reg_2_ (
	.Q(Mfifo_psum_wptr[2]),
	.CK(int_clk),
	.D(Mfifo_psum_M_wptr_wgraynext[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_wptr_wptr_reg_3_ (
	.Q(Mfifo_psum_wptr[3]),
	.CK(int_clk),
	.D(Mfifo_psum_M_wptr_wgraynext[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_wptr_wptr_reg_4_ (
	.Q(Mfifo_psum_wptr[4]),
	.CK(int_clk),
	.D(Mfifo_psum_M_wptr_wbinnext[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_wptr_wbin_reg_0_ (
	.Q(Mfifo_psum_waddr[0]),
	.CK(int_clk),
	.D(Mfifo_psum_M_wptr_wbinnext[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_wptr_wbin_reg_1_ (
	.Q(Mfifo_psum_waddr[1]),
	.CK(int_clk),
	.D(Mfifo_psum_M_wptr_wbinnext[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_wptr_wbin_reg_2_ (
	.Q(Mfifo_psum_waddr[2]),
	.CK(int_clk),
	.D(Mfifo_psum_M_wptr_wbinnext[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_wptr_wbin_reg_3_ (
	.Q(Mfifo_psum_waddr[3]),
	.CK(int_clk),
	.D(Mfifo_psum_M_wptr_wbinnext[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_wptr_wptr_reg_0_ (
	.Q(Mfifo_xin_wptr[0]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_wptr_wgraynext[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_wptr_wptr_reg_1_ (
	.Q(Mfifo_xin_wptr[1]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_wptr_wgraynext[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_wptr_wptr_reg_2_ (
	.Q(Mfifo_xin_wptr[2]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_wptr_wgraynext[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_wptr_wptr_reg_3_ (
	.Q(Mfifo_xin_wptr[3]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_wptr_wgraynext[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_wptr_wptr_reg_4_ (
	.Q(Mfifo_xin_wptr[4]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_wptr_wbinnext[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_wptr_wbin_reg_0_ (
	.Q(Mfifo_xin_waddr[0]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_wptr_wbinnext[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_wptr_wbin_reg_1_ (
	.Q(Mfifo_xin_waddr[1]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_wptr_wbinnext[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_wptr_wbin_reg_2_ (
	.Q(Mfifo_xin_waddr[2]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_wptr_wbinnext[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_wptr_wbin_reg_3_ (
	.Q(Mfifo_xin_waddr[3]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_wptr_wbinnext[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq3_reg_0_ (
	.Q(Mfifo_psum_M_r2w_wq3[0]),
	.CK(int_clk),
	.D(Mfifo_psum_rptr[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq2_reg_0_ (
	.Q(Mfifo_psum_M_r2w_wq2[0]),
	.CK(int_clk),
	.D(Mfifo_psum_M_r2w_wq3[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq2_rptr_reg_0_ (
	.Q(Mfifo_psum_wq2_rptr[0]),
	.CK(int_clk),
	.D(Mfifo_psum_M_r2w_wq2[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq3_reg_1_ (
	.Q(Mfifo_psum_M_r2w_wq3[1]),
	.CK(int_clk),
	.D(Mfifo_psum_rptr[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq2_reg_1_ (
	.Q(Mfifo_psum_M_r2w_wq2[1]),
	.CK(int_clk),
	.D(Mfifo_psum_M_r2w_wq3[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq2_rptr_reg_1_ (
	.Q(Mfifo_psum_wq2_rptr[1]),
	.CK(int_clk),
	.D(Mfifo_psum_M_r2w_wq2[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq3_reg_2_ (
	.Q(Mfifo_psum_M_r2w_wq3[2]),
	.CK(int_clk),
	.D(Mfifo_psum_rptr[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq2_reg_2_ (
	.Q(Mfifo_psum_M_r2w_wq2[2]),
	.CK(int_clk),
	.D(Mfifo_psum_M_r2w_wq3[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq2_rptr_reg_2_ (
	.Q(Mfifo_psum_wq2_rptr[2]),
	.CK(int_clk),
	.D(Mfifo_psum_M_r2w_wq2[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq3_reg_3_ (
	.Q(Mfifo_psum_M_r2w_wq3[3]),
	.CK(int_clk),
	.D(Mfifo_psum_rptr[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq2_reg_3_ (
	.Q(Mfifo_psum_M_r2w_wq2[3]),
	.CK(int_clk),
	.D(Mfifo_psum_M_r2w_wq3[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq2_rptr_reg_3_ (
	.Q(Mfifo_psum_wq2_rptr[3]),
	.CK(int_clk),
	.D(Mfifo_psum_M_r2w_wq2[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq3_reg_4_ (
	.Q(Mfifo_psum_M_r2w_wq3[4]),
	.CK(int_clk),
	.D(Mfifo_psum_rptr[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq2_reg_4_ (
	.Q(Mfifo_psum_M_r2w_wq2[4]),
	.CK(int_clk),
	.D(Mfifo_psum_M_r2w_wq3[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_r2w_wq2_rptr_reg_4_ (
	.Q(Mfifo_psum_wq2_rptr[4]),
	.CK(int_clk),
	.D(Mfifo_psum_M_r2w_wq2[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_wptr_wfull_reg (
	.Q(psum_wfull),
	.CK(int_clk),
	.D(Mfifo_psum_M_wptr_wfull_val),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq3_reg_0_ (
	.Q(Mfifo_xin_M_r2w_wq3[0]),
	.CK(ext_clk),
	.D(Mfifo_xin_rptr[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq2_reg_0_ (
	.Q(Mfifo_xin_M_r2w_wq2[0]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_r2w_wq3[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq2_rptr_reg_0_ (
	.Q(Mfifo_xin_wq2_rptr[0]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_r2w_wq2[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq3_reg_1_ (
	.Q(Mfifo_xin_M_r2w_wq3[1]),
	.CK(ext_clk),
	.D(Mfifo_xin_rptr[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq2_reg_1_ (
	.Q(Mfifo_xin_M_r2w_wq2[1]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_r2w_wq3[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq2_rptr_reg_1_ (
	.Q(Mfifo_xin_wq2_rptr[1]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_r2w_wq2[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq3_reg_2_ (
	.Q(Mfifo_xin_M_r2w_wq3[2]),
	.CK(ext_clk),
	.D(Mfifo_xin_rptr[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq2_reg_2_ (
	.Q(Mfifo_xin_M_r2w_wq2[2]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_r2w_wq3[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq2_rptr_reg_2_ (
	.Q(Mfifo_xin_wq2_rptr[2]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_r2w_wq2[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq3_reg_3_ (
	.Q(Mfifo_xin_M_r2w_wq3[3]),
	.CK(ext_clk),
	.D(Mfifo_xin_rptr[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq2_reg_3_ (
	.Q(Mfifo_xin_M_r2w_wq2[3]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_r2w_wq3[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq2_rptr_reg_3_ (
	.Q(Mfifo_xin_wq2_rptr[3]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_r2w_wq2[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq3_reg_4_ (
	.Q(Mfifo_xin_M_r2w_wq3[4]),
	.CK(ext_clk),
	.D(Mfifo_xin_rptr[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq2_reg_4_ (
	.Q(Mfifo_xin_M_r2w_wq2[4]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_r2w_wq3[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_r2w_wq2_rptr_reg_4_ (
	.Q(Mfifo_xin_wq2_rptr[4]),
	.CK(ext_clk),
	.D(Mfifo_xin_M_r2w_wq2[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_wptr_wfull_reg (
	.Q(n3846),
	.CK(ext_clk),
	.D(Mfifo_xin_M_wptr_wfull_val),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq3_reg_0_ (
	.Q(Mfifo_psum_M_w2r_rq3[0]),
	.CK(ext_clk),
	.D(Mfifo_psum_wptr[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq2_reg_0_ (
	.Q(Mfifo_psum_M_w2r_rq2[0]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_w2r_rq3[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq2_wptr_reg_0_ (
	.Q(Mfifo_psum_rq2_wptr[0]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_w2r_rq2[0]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq3_reg_1_ (
	.Q(Mfifo_psum_M_w2r_rq3[1]),
	.CK(ext_clk),
	.D(Mfifo_psum_wptr[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq2_reg_1_ (
	.Q(Mfifo_psum_M_w2r_rq2[1]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_w2r_rq3[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq2_wptr_reg_1_ (
	.Q(Mfifo_psum_rq2_wptr[1]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_w2r_rq2[1]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq3_reg_2_ (
	.Q(Mfifo_psum_M_w2r_rq3[2]),
	.CK(ext_clk),
	.D(Mfifo_psum_wptr[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq2_reg_2_ (
	.Q(Mfifo_psum_M_w2r_rq2[2]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_w2r_rq3[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq2_wptr_reg_2_ (
	.Q(Mfifo_psum_rq2_wptr[2]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_w2r_rq2[2]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq3_reg_3_ (
	.Q(Mfifo_psum_M_w2r_rq3[3]),
	.CK(ext_clk),
	.D(Mfifo_psum_wptr[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq2_reg_3_ (
	.Q(Mfifo_psum_M_w2r_rq2[3]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_w2r_rq3[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq2_wptr_reg_3_ (
	.Q(Mfifo_psum_rq2_wptr[3]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_w2r_rq2[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq3_reg_4_ (
	.Q(Mfifo_psum_M_w2r_rq3[4]),
	.CK(ext_clk),
	.D(Mfifo_psum_wptr[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq2_reg_4_ (
	.Q(Mfifo_psum_M_w2r_rq2[4]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_w2r_rq3[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_w2r_rq2_wptr_reg_4_ (
	.Q(Mfifo_psum_rq2_wptr[4]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_w2r_rq2[4]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq3_reg_0_ (
	.Q(Mfifo_xin_M_w2r_rq3[0]),
	.CK(int_clk),
	.D(Mfifo_xin_wptr[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq2_reg_0_ (
	.Q(Mfifo_xin_M_w2r_rq2[0]),
	.CK(int_clk),
	.D(Mfifo_xin_M_w2r_rq3[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq2_wptr_reg_0_ (
	.Q(Mfifo_xin_rq2_wptr[0]),
	.CK(int_clk),
	.D(Mfifo_xin_M_w2r_rq2[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq3_reg_1_ (
	.Q(Mfifo_xin_M_w2r_rq3[1]),
	.CK(int_clk),
	.D(Mfifo_xin_wptr[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq2_reg_1_ (
	.Q(Mfifo_xin_M_w2r_rq2[1]),
	.CK(int_clk),
	.D(Mfifo_xin_M_w2r_rq3[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq2_wptr_reg_1_ (
	.Q(Mfifo_xin_rq2_wptr[1]),
	.CK(int_clk),
	.D(Mfifo_xin_M_w2r_rq2[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq3_reg_2_ (
	.Q(Mfifo_xin_M_w2r_rq3[2]),
	.CK(int_clk),
	.D(Mfifo_xin_wptr[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq2_reg_2_ (
	.Q(Mfifo_xin_M_w2r_rq2[2]),
	.CK(int_clk),
	.D(Mfifo_xin_M_w2r_rq3[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq2_wptr_reg_2_ (
	.Q(Mfifo_xin_rq2_wptr[2]),
	.CK(int_clk),
	.D(Mfifo_xin_M_w2r_rq2[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq3_reg_3_ (
	.Q(Mfifo_xin_M_w2r_rq3[3]),
	.CK(int_clk),
	.D(Mfifo_xin_wptr[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq2_reg_3_ (
	.Q(Mfifo_xin_M_w2r_rq2[3]),
	.CK(int_clk),
	.D(Mfifo_xin_M_w2r_rq3[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq2_wptr_reg_3_ (
	.Q(Mfifo_xin_rq2_wptr[3]),
	.CK(int_clk),
	.D(Mfifo_xin_M_w2r_rq2[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq3_reg_4_ (
	.Q(Mfifo_xin_M_w2r_rq3[4]),
	.CK(int_clk),
	.D(Mfifo_xin_wptr[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq2_reg_4_ (
	.Q(Mfifo_xin_M_w2r_rq2[4]),
	.CK(int_clk),
	.D(Mfifo_xin_M_w2r_rq3[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_w2r_rq2_wptr_reg_4_ (
	.Q(Mfifo_xin_rq2_wptr[4]),
	.CK(int_clk),
	.D(Mfifo_xin_M_w2r_rq2[4]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_synsend_sync2_reg (
	.Q(Msyncin_synsend_sync2),
	.CK(int_clk),
	.D(ext_send),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_synsend_sync1_reg (
	.Q(Msyncin_synsend_sync1),
	.CK(int_clk),
	.D(Msyncin_synsend_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_synsend_synced_reg (
	.Q(int_send),
	.CK(int_clk),
	.D(Msyncin_synsend_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_syncomp_sync2_reg (
	.Q(Msyncin_syncomp_sync2),
	.CK(int_clk),
	.D(ext_comp),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_syncomp_sync1_reg (
	.Q(Msyncin_syncomp_sync1),
	.CK(int_clk),
	.D(Msyncin_syncomp_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_syncomp_synced_reg (
	.Q(int_comp),
	.CK(int_clk),
	.D(Msyncin_syncomp_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_synenable_sync2_reg (
	.Q(Msyncin_synenable_sync2),
	.CK(int_clk),
	.D(ext_enable),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_synenable_sync1_reg (
	.Q(Msyncin_synenable_sync1),
	.CK(int_clk),
	.D(Msyncin_synenable_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_synenable_synced_reg (
	.Q(int_enable),
	.CK(int_clk),
	.D(Msyncin_synenable_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_3__synH_sync2_reg (
	.Q(Msyncin_MsynWH_3__synH_sync2),
	.CK(int_clk),
	.D(ext_H[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_3__synH_sync1_reg (
	.Q(Msyncin_MsynWH_3__synH_sync1),
	.CK(int_clk),
	.D(Msyncin_MsynWH_3__synH_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_3__synH_synced_reg (
	.Q(int_H[3]),
	.CK(int_clk),
	.D(Msyncin_MsynWH_3__synH_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_3__synW_sync2_reg (
	.Q(Msyncin_MsynWH_3__synW_sync2),
	.CK(int_clk),
	.D(ext_W[3]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_3__synW_sync1_reg (
	.Q(Msyncin_MsynWH_3__synW_sync1),
	.CK(int_clk),
	.D(Msyncin_MsynWH_3__synW_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_3__synW_synced_reg (
	.Q(int_W[3]),
	.CK(int_clk),
	.D(Msyncin_MsynWH_3__synW_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_2__synH_sync2_reg (
	.Q(Msyncin_MsynWH_2__synH_sync2),
	.CK(int_clk),
	.D(ext_H[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_2__synH_sync1_reg (
	.Q(Msyncin_MsynWH_2__synH_sync1),
	.CK(int_clk),
	.D(Msyncin_MsynWH_2__synH_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_2__synH_synced_reg (
	.Q(int_H[2]),
	.CK(int_clk),
	.D(Msyncin_MsynWH_2__synH_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_2__synW_sync2_reg (
	.Q(Msyncin_MsynWH_2__synW_sync2),
	.CK(int_clk),
	.D(ext_W[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_2__synW_sync1_reg (
	.Q(Msyncin_MsynWH_2__synW_sync1),
	.CK(int_clk),
	.D(Msyncin_MsynWH_2__synW_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_2__synW_synced_reg (
	.Q(int_W[2]),
	.CK(int_clk),
	.D(Msyncin_MsynWH_2__synW_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_1__synH_sync2_reg (
	.Q(Msyncin_MsynWH_1__synH_sync2),
	.CK(int_clk),
	.D(ext_H[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_1__synH_sync1_reg (
	.Q(Msyncin_MsynWH_1__synH_sync1),
	.CK(int_clk),
	.D(Msyncin_MsynWH_1__synH_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_1__synH_synced_reg (
	.Q(int_H[1]),
	.CK(int_clk),
	.D(Msyncin_MsynWH_1__synH_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_1__synW_sync2_reg (
	.Q(Msyncin_MsynWH_1__synW_sync2),
	.CK(int_clk),
	.D(ext_W[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_1__synW_sync1_reg (
	.Q(Msyncin_MsynWH_1__synW_sync1),
	.CK(int_clk),
	.D(Msyncin_MsynWH_1__synW_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_1__synW_synced_reg (
	.Q(int_W[1]),
	.CK(int_clk),
	.D(Msyncin_MsynWH_1__synW_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_0__synH_sync2_reg (
	.Q(Msyncin_MsynWH_0__synH_sync2),
	.CK(int_clk),
	.D(ext_H[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_0__synH_sync1_reg (
	.Q(Msyncin_MsynWH_0__synH_sync1),
	.CK(int_clk),
	.D(Msyncin_MsynWH_0__synH_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_0__synH_synced_reg (
	.Q(int_H[0]),
	.CK(int_clk),
	.D(Msyncin_MsynWH_0__synH_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_0__synW_sync2_reg (
	.Q(Msyncin_MsynWH_0__synW_sync2),
	.CK(int_clk),
	.D(ext_W[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_0__synW_sync1_reg (
	.Q(Msyncin_MsynWH_0__synW_sync1),
	.CK(int_clk),
	.D(Msyncin_MsynWH_0__synW_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_MsynWH_0__synW_synced_reg (
	.Q(int_W[0]),
	.CK(int_clk),
	.D(Msyncin_MsynWH_0__synW_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_1__synky_sync2_reg (
	.Q(Msyncin_Msynkxy_1__synky_sync2),
	.CK(int_clk),
	.D(ext_ky[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_1__synky_sync1_reg (
	.Q(Msyncin_Msynkxy_1__synky_sync1),
	.CK(int_clk),
	.D(Msyncin_Msynkxy_1__synky_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_1__synky_synced_reg (
	.Q(int_ky[1]),
	.CK(int_clk),
	.D(Msyncin_Msynkxy_1__synky_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_1__synkx_sync2_reg (
	.Q(Msyncin_Msynkxy_1__synkx_sync2),
	.CK(int_clk),
	.D(ext_kx[1]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_1__synkx_sync1_reg (
	.Q(Msyncin_Msynkxy_1__synkx_sync1),
	.CK(int_clk),
	.D(Msyncin_Msynkxy_1__synkx_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_1__synkx_synced_reg (
	.Q(int_kx[1]),
	.CK(int_clk),
	.D(Msyncin_Msynkxy_1__synkx_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_0__synky_sync2_reg (
	.Q(Msyncin_Msynkxy_0__synky_sync2),
	.CK(int_clk),
	.D(ext_ky[0]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_0__synky_sync1_reg (
	.Q(Msyncin_Msynkxy_0__synky_sync1),
	.CK(int_clk),
	.D(Msyncin_Msynkxy_0__synky_sync2),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncin_Msynkxy_0__synky_synced_reg (
	.Q(int_ky[0]),
	.CK(int_clk),
	.D(Msyncin_Msynkxy_0__synky_sync1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_ky_reg_0_ (
	.Q(c_ky[0]),
	.CK(int_clk),
	.D(n2385),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_x_cin_reg_0_ (
	.Q(Mcntl_Mcntldata_c_x_cin[0]),
	.CK(int_clk),
	.D(n2081),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntl_current_state_reg_0_ (
	.Q(Mcntl_Mcntl_current_state[0]),
	.CK(int_clk),
	.D(n2395),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_cout_reg_2_ (
	.Q(Mcntl_Mcntldata_c_p_cout[2]),
	.CK(int_clk),
	.D(n2373),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntl_current_state_reg_1_ (
	.Q(Mcntl_Mcntl_current_state[1]),
	.CK(int_clk),
	.D(n2393),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncout_syneread_sync2_reg (
	.Q(Msyncout_syneread_sync2),
	.CK(ext_clk),
	.D(int_end_read),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncout_syneread_sync1_reg (
	.Q(Msyncout_syneread_sync1),
	.CK(ext_clk),
	.D(Msyncout_syneread_sync2),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncout_syneread_synced_reg (
	.Q(ext_end_read),
	.CK(ext_clk),
	.D(Msyncout_syneread_sync1),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntl_current_state_reg_2_ (
	.Q(Mcntl_Mcntl_current_state[2]),
	.CK(int_clk),
	.D(n2394),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncout_synesend_sync2_reg (
	.Q(Msyncout_synesend_sync2),
	.CK(ext_clk),
	.D(int_end_send),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncout_synesend_sync1_reg (
	.Q(Msyncout_synesend_sync1),
	.CK(ext_clk),
	.D(Msyncout_synesend_sync2),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncout_synesend_synced_reg (
	.Q(ext_end_send),
	.CK(ext_clk),
	.D(Msyncout_synesend_sync1),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_cin_reg_0_ (
	.Q(Mcntl_Mcntldata_c_cin[0]),
	.CK(int_clk),
	.D(n2377),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_cin_reg_1_ (
	.Q(Mcntl_Mcntldata_c_cin[1]),
	.CK(int_clk),
	.D(n2378),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_cout_reg_0_ (
	.Q(c_cout[0]),
	.CK(int_clk),
	.D(n2383),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_cout_reg_1_ (
	.Q(c_cout[1]),
	.CK(int_clk),
	.D(n2382),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_cout_reg_2_ (
	.Q(c_cout[2]),
	.CK(int_clk),
	.D(n2381),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_cout_reg_3_ (
	.Q(c_cout[3]),
	.CK(int_clk),
	.D(n2380),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_kx_reg_0_ (
	.Q(c_kx[0]),
	.CK(int_clk),
	.D(n2379),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_ky_reg_1_ (
	.Q(c_ky[1]),
	.CK(int_clk),
	.D(n2386),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_kx_reg_1_ (
	.Q(c_kx[1]),
	.CK(int_clk),
	.D(n2392),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_flag_reg (
	.Q(Mcntl_flag),
	.CK(int_clk),
	.D(n2376),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_count_reg_1_ (
	.Q(Mcntl_Mcntldata_count[1]),
	.CK(int_clk),
	.D(n2390),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_count_reg_0_ (
	.Q(Mcntl_Mcntldata_count[0]),
	.CK(int_clk),
	.D(n2391),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_count_k_reg_2_ (
	.Q(count_k[2]),
	.CK(int_clk),
	.D(n2387),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_count_k_reg_0_ (
	.Q(count_k[0]),
	.CK(int_clk),
	.D(n2388),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_count_k_reg_1_ (
	.Q(count_k[1]),
	.CK(int_clk),
	.D(n2389),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_wd4_reg_1_ (
	.Q(Mcntl_Mcntldata_c_p_wd4[1]),
	.CK(int_clk),
	.D(n2364),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_wd4_reg_0_ (
	.Q(Mcntl_Mcntldata_c_p_wd4[0]),
	.CK(int_clk),
	.D(n2365),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_comp_psum_reg (
	.Q(Mcntl_Mcntldata_comp_psum),
	.CK(int_clk),
	.D(n2079),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncout_synepsum_sync2_reg (
	.Q(Msyncout_synepsum_sync2),
	.CK(ext_clk),
	.D(int_end_comp),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncout_synepsum_sync1_reg (
	.Q(Msyncout_synepsum_sync1),
	.CK(ext_clk),
	.D(Msyncout_synepsum_sync2),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Msyncout_synepsum_synced_reg (
	.Q(ext_end_comp),
	.CK(ext_clk),
	.D(Msyncout_synepsum_sync1),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_cout_reg_1_ (
	.Q(Mcntl_Mcntldata_c_p_cout[1]),
	.CK(int_clk),
	.D(n2375),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_W_reg_0_ (
	.Q(sel_reg[0]),
	.CK(int_clk),
	.D(n2370),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_W_reg_1_ (
	.Q(sel_reg[1]),
	.CK(int_clk),
	.D(n2372),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_W_reg_2_ (
	.Q(Mcntl_Mcntldata_c_p_W[2]),
	.CK(int_clk),
	.D(n2371),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_W_reg_3_ (
	.Q(Mcntl_Mcntldata_c_p_W[3]),
	.CK(int_clk),
	.D(n2384),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_H_reg_3_ (
	.Q(Mcntl_Mcntldata_c_p_H[3]),
	.CK(int_clk),
	.D(n2366),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_H_reg_0_ (
	.Q(Mcntl_Mcntldata_c_p_H[0]),
	.CK(int_clk),
	.D(n2369),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_H_reg_1_ (
	.Q(Mcntl_Mcntldata_c_p_H[1]),
	.CK(int_clk),
	.D(n2368),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_H_reg_2_ (
	.Q(Mcntl_Mcntldata_c_p_H[2]),
	.CK(int_clk),
	.D(n2367),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_cin_reg_0_ (
	.Q(Mcntl_Mcntldata_c_p_cin[0]),
	.CK(int_clk),
	.D(n2363),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_p_cin_reg_1_ (
	.Q(Mcntl_Mcntldata_c_p_cin[1]),
	.CK(int_clk),
	.D(n2362),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_W_r4_reg_0_ (
	.Q(Mcntl_Mcntldata_c_W_r4[0]),
	.CK(int_clk),
	.D(n2080),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_W_d4_reg_0_ (
	.Q(Mcntl_Mcntldata_c_W_d4[0]),
	.CK(int_clk),
	.D(n2083),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_W_d4_reg_1_ (
	.Q(Mcntl_Mcntldata_c_W_d4[1]),
	.CK(int_clk),
	.D(n2089),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 R_21128 (
	.Q(Mcntl_Mcntldata_c_x_H[0]),
	.CK(int_clk),
	.D(n2084),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_x_H_reg_3_ (
	.Q(Mcntl_Mcntldata_c_x_H[3]),
	.CK(int_clk),
	.D(n2087),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_x_H_reg_2_ (
	.Q(Mcntl_Mcntldata_c_x_H[2]),
	.CK(int_clk),
	.D(n2086),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 R_21129 (
	.Q(Mcntl_Mcntldata_c_x_H[1]),
	.CK(int_clk),
	.D(n2085),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_x_cin_reg_1_ (
	.Q(Mcntl_Mcntldata_c_x_cin[1]),
	.CK(int_clk),
	.D(n2082),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_c_W_r4_reg_1_ (
	.Q(Mcntl_Mcntldata_c_W_r4[1]),
	.CK(int_clk),
	.D(n2088),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_addr_reg_1_ (
	.Q(x_addr[1]),
	.CK(int_clk),
	.D(n2072),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_addr_reg_0_ (
	.Q(x_addr[0]),
	.CK(int_clk),
	.D(n2071),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_addr_reg_2_ (
	.Q(x_addr[2]),
	.CK(int_clk),
	.D(n2070),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_addr_reg_3_ (
	.Q(x_addr[3]),
	.CK(int_clk),
	.D(n2069),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_addr_reg_4_ (
	.Q(x_addr[4]),
	.CK(int_clk),
	.D(n2068),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_addr_reg_5_ (
	.Q(x_addr[5]),
	.CK(int_clk),
	.D(n2067),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_addr_reg_6_ (
	.Q(x_addr[6]),
	.CK(int_clk),
	.D(n3832),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntl_Mwenc_qout_r_reg_0_ (
	.Q(wen_coe),
	.CK(int_clk),
	.D(Mfifo_coe_M_rptr_N1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntl_Mwenx_qout_r_reg_0_ (
	.Q(wen_x),
	.CK(int_clk),
	.D(Mfifo_xin_M_rptr_N1),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX1AR9 Mfifo_coe_M_ffmem_rdata_reg_1_ (
	.Q(int_coe[1]),
	.CK(int_clk),
	.D(n2233), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX1AR9 Mfifo_coe_M_ffmem_rdata_reg_3_ (
	.Q(int_coe[3]),
	.CK(int_clk),
	.D(n2231), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX1AR9 Mfifo_coe_M_ffmem_rdata_reg_4_ (
	.Q(int_coe[4]),
	.CK(int_clk),
	.D(n2230), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX1AR9 Mfifo_coe_M_ffmem_rdata_reg_7_ (
	.Q(int_coe[7]),
	.CK(int_clk),
	.D(n2227), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX1AR9 Mfifo_coe_M_ffmem_rdata_reg_0_ (
	.Q(int_coe[0]),
	.CK(int_clk),
	.D(n2226), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFSBQX05AR9 Mfifo_coe_M_rptr_rempty_reg (
	.Q(coe_rempty),
	.CK(int_clk),
	.D(Mfifo_coe_M_rptr_rempty_val),
	.SB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFSBQX05AR9 Mfifo_psum_M_rptr_rempty_reg (
	.Q(n3847),
	.CK(ext_clk),
	.D(Mfifo_psum_M_rptr_rempty_val),
	.SB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFSBQX05AR9 Mfifo_xin_M_rptr_rempty_reg (
	.Q(xin_rempty),
	.CK(int_clk),
	.D(Mfifo_xin_M_rptr_rempty_val),
	.SB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_kx_reg_reg_1_ (
	.Q(Mcntl_Mcntldata_kx_reg[1]),
	.CK(int_clk),
	.D(n1393),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_ky_reg_reg_0_ (
	.Q(Mcntl_Mcntldata_ky_reg[0]),
	.CK(int_clk),
	.D(n1392),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_ky_reg_reg_1_ (
	.Q(Mcntl_Mcntldata_ky_reg[1]),
	.CK(int_clk),
	.D(n1391),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_W_reg_reg_0_ (
	.Q(Mcntl_Mcntldata_x_W_reg[0]),
	.CK(int_clk),
	.D(n1390),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_W_reg_reg_1_ (
	.Q(Mcntl_Mcntldata_x_W_reg[1]),
	.CK(int_clk),
	.D(n1389),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_W_reg_reg_2_ (
	.Q(Mcntl_Mcntldata_x_W_reg[2]),
	.CK(int_clk),
	.D(n1388),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_W_reg_reg_3_ (
	.Q(Mcntl_Mcntldata_x_W_reg[3]),
	.CK(int_clk),
	.D(n1387),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_H_reg_reg_0_ (
	.Q(Mcntl_Mcntldata_x_H_reg[0]),
	.CK(int_clk),
	.D(n1386),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_H_reg_reg_1_ (
	.Q(Mcntl_Mcntldata_x_H_reg[1]),
	.CK(int_clk),
	.D(n1385),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_H_reg_reg_2_ (
	.Q(Mcntl_Mcntldata_x_H_reg[2]),
	.CK(int_clk),
	.D(n1384),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_x_H_reg_reg_3_ (
	.Q(Mcntl_Mcntldata_x_H_reg[3]),
	.CK(int_clk),
	.D(n1383),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_kx_reg_reg_0_ (
	.Q(Mcntl_Mcntldata_kx_reg[0]),
	.CK(int_clk),
	.D(n1382),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_0 MRegpsum_Mpsumreg4_4 (
	.dataout(psum4_reg4),
	.datain(psum4_o4),
	.addr({ n3843,
		psum_addr[4],
		n3834,
		n3840,
		n3837,
		n3838 }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_1 MRegpsum_Mpsumreg4_3 (
	.dataout(psum4_reg3),
	.datain(psum4_o3),
	.addr({ n3843,
		psum_addr[4],
		n3834,
		n3831,
		n3836,
		psum_addr[0] }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_2 MRegpsum_Mpsumreg4_2 (
	.dataout(psum4_reg2),
	.datain(psum4_o2),
	.addr({ n3843,
		psum_addr[4],
		n3835,
		n3831,
		n3836,
		n3838 }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_3 MRegpsum_Mpsumreg4_1 (
	.dataout(psum4_reg1),
	.datain(psum4_o1),
	.addr({ n3843,
		psum_addr[4],
		n3835,
		n3831,
		psum_addr[1],
		psum_addr[0] }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_4 MRegpsum_Mpsumreg3_4 (
	.dataout(psum3_reg4),
	.datain(psum3_o4),
	.addr({ n3843,
		psum_addr[4],
		n3834,
		n3840,
		psum_addr[1],
		psum_addr[0] }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_5 MRegpsum_Mpsumreg3_3 (
	.dataout(psum3_reg3),
	.datain(psum3_o3),
	.addr({ n3843,
		psum_addr[4],
		n3834,
		n3841,
		n3837,
		psum_addr[0] }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_6 MRegpsum_Mpsumreg3_2 (
	.dataout(psum3_reg2),
	.datain(psum3_o2),
	.addr({ n3843,
		psum_addr[4],
		n3834,
		n2076,
		n3836,
		psum_addr[0] }),
	.write(n2413),
	.clk(int_clk),
	.IN0(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_7 MRegpsum_Mpsumreg3_1 (
	.dataout(psum3_reg1),
	.datain(psum3_o1),
	.addr({ n3843,
		psum_addr[4],
		n3834,
		n3841,
		psum_addr[1],
		psum_addr[0] }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_8 MRegpsum_Mpsumreg2_4 (
	.dataout(psum2_reg4),
	.datain(psum2_o4),
	.addr({ n3843,
		psum_addr[4],
		n3834,
		n3830,
		n3837,
		n3838 }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_9 MRegpsum_Mpsumreg2_3 (
	.dataout(psum2_reg3),
	.datain(psum2_o3),
	.addr({ n3843,
		psum_addr[4],
		n3834,
		n3841,
		n3836,
		psum_addr[0] }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_10 MRegpsum_Mpsumreg2_2 (
	.dataout(psum2_reg2),
	.datain(psum2_o2),
	.addr({ n3843,
		psum_addr[4],
		n3834,
		n3830,
		n3836,
		psum_addr[0] }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_11 MRegpsum_Mpsumreg2_1 (
	.dataout(psum2_reg1),
	.datain(psum2_o1),
	.addr({ n3843,
		psum_addr[4],
		n3834,
		n3841,
		n3836,
		psum_addr[0] }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_12 MRegpsum_Mpsumreg1_4 (
	.dataout(psum1_reg4),
	.datain(psum1_o4),
	.addr({ psum_addr[5],
		psum_addr[4],
		n3834,
		n3830,
		psum_addr[1],
		n2077 }),
	.write(n2413),
	.clk(int_clk),
	.IN0(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_13 MRegpsum_Mpsumreg1_3 (
	.dataout(psum1_reg3),
	.datain(psum1_o3),
	.addr({ psum_addr[5],
		psum_addr[4],
		n3834,
		n3841,
		n3836,
		psum_addr[0] }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_14 MRegpsum_Mpsumreg1_2 (
	.dataout(psum1_reg2),
	.datain(psum1_o2),
	.addr({ psum_addr[5],
		psum_addr[4],
		n3834,
		n3841,
		n3836,
		n3838 }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   Reg_psum_file_mini_15 MRegpsum_Mpsumreg1_1 (
	.dataout(psum1_reg1),
	.datain(psum1_o1),
	.addr({ psum_addr[5],
		psum_addr[4],
		n3834,
		n3831,
		psum_addr[1],
		psum_addr[0] }),
	.write(n2413),
	.clk(int_clk), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 DP_OP_1205J5_125_5849_U8 (
	.CO(DP_OP_1205J5_125_5849_n7),
	.S(C174_DATA2_0),
	.CI(DP_OP_1205J5_125_5849_n15),
	.I1(C2_Z_0),
	.I2(x_addr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 DP_OP_1205J5_125_5849_U7 (
	.CO(DP_OP_1205J5_125_5849_n6),
	.S(C174_DATA2_1),
	.CI(DP_OP_1205J5_125_5849_n7),
	.I1(x_addr[1]),
	.I2(DP_OP_1205J5_125_5849_n14), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 DP_OP_1205J5_125_5849_U6 (
	.CO(DP_OP_1205J5_125_5849_n5),
	.S(C174_DATA2_2),
	.CI(DP_OP_1205J5_125_5849_n6),
	.I1(x_addr[2]),
	.I2(DP_OP_1205J5_125_5849_n13), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 DP_OP_1205J5_125_5849_U5 (
	.CO(DP_OP_1205J5_125_5849_n4),
	.S(C174_DATA2_3),
	.CI(DP_OP_1205J5_125_5849_n5),
	.I1(x_addr[3]),
	.I2(DP_OP_1205J5_125_5849_n12), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 DP_OP_1205J5_125_5849_U4 (
	.CO(DP_OP_1205J5_125_5849_n3),
	.S(C174_DATA2_4),
	.CI(DP_OP_1205J5_125_5849_n4),
	.I1(x_addr[4]),
	.I2(C2_Z_0), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 DP_OP_1205J5_125_5849_U3 (
	.CO(DP_OP_1205J5_125_5849_n2),
	.S(C174_DATA2_5),
	.CI(DP_OP_1205J5_125_5849_n3),
	.I1(x_addr[5]),
	.I2(C2_Z_0), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 DP_OP_1207J5_130_8771_U5 (
	.CO(DP_OP_1207J5_130_8771_n4),
	.S(C175_DATA2_2),
	.CI(n3833),
	.I1(n3841),
	.I2(Mcntl_Mcntldata_N453), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_psum_M_rptr_rbin_reg_3_ (
	.Q(Mfifo_psum_raddr[3]),
	.CK(ext_clk),
	.D(Mfifo_psum_M_rptr_rbinnext[3]),
	.RB(ext_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mfifo_xin_M_rptr_rbin_reg_2_ (
	.Q(Mfifo_xin_raddr[2]),
	.CK(int_clk),
	.D(Mfifo_xin_M_rptr_rbinnext[2]),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX8K1AR9 Mcntl_Mcntldata_psum_addr_reg_4_ (
	.Q(psum_addr[4]),
	.CK(int_clk),
	.D(n2074),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX4K1AR9 R_21189 (
	.Q(n3840),
	.CK(int_clk),
	.D(n2076),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_21_ (
	.Q(ext_psum2[0]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N96),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_22_ (
	.Q(ext_psum2[1]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N95),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_23_ (
	.Q(ext_psum2[2]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N94),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_24_ (
	.Q(ext_psum2[3]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N93),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_25_ (
	.Q(ext_psum2[4]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N92),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_26_ (
	.Q(ext_psum2[5]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N91),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_27_ (
	.Q(ext_psum2[6]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N90),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_28_ (
	.Q(ext_psum2[7]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N89),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_29_ (
	.Q(ext_psum2[8]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N88),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_30_ (
	.Q(ext_psum2[9]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N87),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_31_ (
	.Q(ext_psum2[10]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N86),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_32_ (
	.Q(ext_psum2[11]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N85),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_33_ (
	.Q(ext_psum2[12]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N84),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_34_ (
	.Q(ext_psum2[13]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N83),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_35_ (
	.Q(ext_psum2[14]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N82),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_36_ (
	.Q(ext_psum2[15]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N81),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_37_ (
	.Q(ext_psum2[16]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N80),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_38_ (
	.Q(ext_psum2[17]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N79),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_39_ (
	.Q(ext_psum2[18]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N78),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_40_ (
	.Q(ext_psum2[19]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N77),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_41_ (
	.Q(ext_psum2[20]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N76),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_0_ (
	.Q(ext_psum1[0]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N117),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_1_ (
	.Q(ext_psum1[1]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N116),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_2_ (
	.Q(ext_psum1[2]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N115),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_3_ (
	.Q(ext_psum1[3]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N114),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_4_ (
	.Q(ext_psum1[4]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N113),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_5_ (
	.Q(ext_psum1[5]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N112),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_6_ (
	.Q(ext_psum1[6]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N111),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_7_ (
	.Q(ext_psum1[7]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N110),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_8_ (
	.Q(ext_psum1[8]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N109),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_9_ (
	.Q(ext_psum1[9]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N108),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_10_ (
	.Q(ext_psum1[10]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N107),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_11_ (
	.Q(ext_psum1[11]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N106),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_12_ (
	.Q(ext_psum1[12]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N105),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_13_ (
	.Q(ext_psum1[13]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N104),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_14_ (
	.Q(ext_psum1[14]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N103),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_15_ (
	.Q(ext_psum1[15]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N102),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_16_ (
	.Q(ext_psum1[16]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N101),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_17_ (
	.Q(ext_psum1[17]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N100),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_18_ (
	.Q(ext_psum1[18]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N99),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_19_ (
	.Q(ext_psum1[19]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N98),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFCNLDQX05AR9 Mfifo_psum_M_ffmem_rdata_reg_20_ (
	.Q(ext_psum1[20]),
	.CK(ext_clk),
	.CN(1'b1),
	.D(Mfifo_psum_M_ffmem_N97),
	.LD(n3842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_15__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_15__6_),
	.CK(ext_clk),
	.D(n2359), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_11__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_11__7_),
	.CK(ext_clk),
	.D(n2328), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_14__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_14__0_),
	.CK(ext_clk),
	.D(n2353), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_12__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_12__1_),
	.CK(ext_clk),
	.D(n2330), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_8__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_8__2_),
	.CK(ext_clk),
	.D(n2299), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_5__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_5__3_),
	.CK(ext_clk),
	.D(n2276), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_1__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_1__4_),
	.CK(ext_clk),
	.D(n2245), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_4__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_4__5_),
	.CK(ext_clk),
	.D(n2270), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_0__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_0__6_),
	.CK(ext_clk),
	.D(n2239), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_13__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_13__7_),
	.CK(ext_clk),
	.D(n2208), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_9__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_9__0_),
	.CK(ext_clk),
	.D(n2177), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_14__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_14__1_),
	.CK(ext_clk),
	.D(n2210), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_10__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_10__2_),
	.CK(ext_clk),
	.D(n2179), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_7__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_7__3_),
	.CK(ext_clk),
	.D(n2156), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_3__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_3__4_),
	.CK(ext_clk),
	.D(n2125), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_6__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_6__5_),
	.CK(ext_clk),
	.D(n2150), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_2__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_2__6_),
	.CK(ext_clk),
	.D(n2119), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__21_),
	.CK(int_clk),
	.D(n2065), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__21_),
	.CK(int_clk),
	.D(n2050), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__22_),
	.CK(int_clk),
	.D(n2035), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__23_),
	.CK(int_clk),
	.D(n2020), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__24_),
	.CK(int_clk),
	.D(n2005), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__25_),
	.CK(int_clk),
	.D(n1990), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__26_),
	.CK(int_clk),
	.D(n1975), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__27_),
	.CK(int_clk),
	.D(n1960), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__28_),
	.CK(int_clk),
	.D(n1945), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__29_),
	.CK(int_clk),
	.D(n1930), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__30_),
	.CK(int_clk),
	.D(n1915), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__31_),
	.CK(int_clk),
	.D(n1900), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__32_),
	.CK(int_clk),
	.D(n1885), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__33_),
	.CK(int_clk),
	.D(n1870), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__34_),
	.CK(int_clk),
	.D(n1855), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__35_),
	.CK(int_clk),
	.D(n1840), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__36_),
	.CK(int_clk),
	.D(n1825), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__36_),
	.CK(int_clk),
	.D(n1810), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__37_),
	.CK(int_clk),
	.D(n1795), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__38_),
	.CK(int_clk),
	.D(n1780), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__39_),
	.CK(int_clk),
	.D(n1765), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__40_),
	.CK(int_clk),
	.D(n1750), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__41_),
	.CK(int_clk),
	.D(n1735), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__0_),
	.CK(int_clk),
	.D(n1720), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__1_),
	.CK(int_clk),
	.D(n1705), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__2_),
	.CK(int_clk),
	.D(n1690), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__3_),
	.CK(int_clk),
	.D(n1675), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__4_),
	.CK(int_clk),
	.D(n1660), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__5_),
	.CK(int_clk),
	.D(n1645), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__6_),
	.CK(int_clk),
	.D(n1630), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__7_),
	.CK(int_clk),
	.D(n1615), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__8_),
	.CK(int_clk),
	.D(n1600), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__9_),
	.CK(int_clk),
	.D(n1585), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__9_),
	.CK(int_clk),
	.D(n1570), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__10_),
	.CK(int_clk),
	.D(n1555), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__11_),
	.CK(int_clk),
	.D(n1540), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__12_),
	.CK(int_clk),
	.D(n1525), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__13_),
	.CK(int_clk),
	.D(n1510), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__14_),
	.CK(int_clk),
	.D(n1495), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__15_),
	.CK(int_clk),
	.D(n1480), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__16_),
	.CK(int_clk),
	.D(n1465), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__17_),
	.CK(int_clk),
	.D(n1450), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__18_),
	.CK(int_clk),
	.D(n1435), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__19_),
	.CK(int_clk),
	.D(n1420), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__20_),
	.CK(int_clk),
	.D(n1405), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__20_),
	.CK(int_clk),
	.D(n1394), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 R_20584 (
	.Q(psum_addr[5]),
	.CK(int_clk),
	.D(n2073),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_15__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_15__0_),
	.CK(ext_clk),
	.D(n2361), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_15__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_15__7_),
	.CK(ext_clk),
	.D(n2360), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_15__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_15__5_),
	.CK(ext_clk),
	.D(n2358), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_15__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_15__4_),
	.CK(ext_clk),
	.D(n2357), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_15__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_15__3_),
	.CK(ext_clk),
	.D(n2356), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_15__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_15__2_),
	.CK(ext_clk),
	.D(n2355), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_15__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_15__1_),
	.CK(ext_clk),
	.D(n2354), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_13__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_13__0_),
	.CK(ext_clk),
	.D(n2345), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_13__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_13__7_),
	.CK(ext_clk),
	.D(n2344), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_13__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_13__6_),
	.CK(ext_clk),
	.D(n2343), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_13__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_13__5_),
	.CK(ext_clk),
	.D(n2342), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_13__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_13__4_),
	.CK(ext_clk),
	.D(n2341), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_13__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_13__3_),
	.CK(ext_clk),
	.D(n2340), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_13__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_13__2_),
	.CK(ext_clk),
	.D(n2339), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_13__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_13__1_),
	.CK(ext_clk),
	.D(n2338), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_11__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_11__0_),
	.CK(ext_clk),
	.D(n2329), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_11__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_11__6_),
	.CK(ext_clk),
	.D(n2327), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_11__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_11__5_),
	.CK(ext_clk),
	.D(n2326), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_11__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_11__4_),
	.CK(ext_clk),
	.D(n2325), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_11__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_11__3_),
	.CK(ext_clk),
	.D(n2324), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_11__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_11__2_),
	.CK(ext_clk),
	.D(n2323), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_11__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_11__1_),
	.CK(ext_clk),
	.D(n2322), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_9__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_9__0_),
	.CK(ext_clk),
	.D(n2313), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_9__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_9__7_),
	.CK(ext_clk),
	.D(n2312), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_9__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_9__6_),
	.CK(ext_clk),
	.D(n2311), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_9__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_9__5_),
	.CK(ext_clk),
	.D(n2310), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_9__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_9__4_),
	.CK(ext_clk),
	.D(n2309), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_9__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_9__3_),
	.CK(ext_clk),
	.D(n2308), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_9__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_9__2_),
	.CK(ext_clk),
	.D(n2307), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_9__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_9__1_),
	.CK(ext_clk),
	.D(n2306), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_14__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_14__7_),
	.CK(ext_clk),
	.D(n2352), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_14__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_14__6_),
	.CK(ext_clk),
	.D(n2351), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_14__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_14__5_),
	.CK(ext_clk),
	.D(n2350), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_14__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_14__4_),
	.CK(ext_clk),
	.D(n2349), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_14__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_14__3_),
	.CK(ext_clk),
	.D(n2348), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_14__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_14__2_),
	.CK(ext_clk),
	.D(n2347), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_14__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_14__1_),
	.CK(ext_clk),
	.D(n2346), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_12__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_12__0_),
	.CK(ext_clk),
	.D(n2337), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_12__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_12__7_),
	.CK(ext_clk),
	.D(n2336), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_12__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_12__6_),
	.CK(ext_clk),
	.D(n2335), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_12__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_12__5_),
	.CK(ext_clk),
	.D(n2334), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_12__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_12__4_),
	.CK(ext_clk),
	.D(n2333), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_12__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_12__3_),
	.CK(ext_clk),
	.D(n2332), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_12__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_12__2_),
	.CK(ext_clk),
	.D(n2331), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_10__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_10__0_),
	.CK(ext_clk),
	.D(n2321), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_10__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_10__7_),
	.CK(ext_clk),
	.D(n2320), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_10__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_10__6_),
	.CK(ext_clk),
	.D(n2319), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_10__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_10__5_),
	.CK(ext_clk),
	.D(n2318), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_10__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_10__4_),
	.CK(ext_clk),
	.D(n2317), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_10__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_10__3_),
	.CK(ext_clk),
	.D(n2316), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_10__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_10__2_),
	.CK(ext_clk),
	.D(n2315), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_10__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_10__1_),
	.CK(ext_clk),
	.D(n2314), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_8__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_8__0_),
	.CK(ext_clk),
	.D(n2305), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_8__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_8__7_),
	.CK(ext_clk),
	.D(n2304), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_8__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_8__6_),
	.CK(ext_clk),
	.D(n2303), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_8__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_8__5_),
	.CK(ext_clk),
	.D(n2302), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_8__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_8__4_),
	.CK(ext_clk),
	.D(n2301), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_8__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_8__3_),
	.CK(ext_clk),
	.D(n2300), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_8__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_8__1_),
	.CK(ext_clk),
	.D(n2298), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_7__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_7__0_),
	.CK(ext_clk),
	.D(n2297), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_7__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_7__7_),
	.CK(ext_clk),
	.D(n2296), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_7__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_7__6_),
	.CK(ext_clk),
	.D(n2295), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_7__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_7__5_),
	.CK(ext_clk),
	.D(n2294), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_7__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_7__4_),
	.CK(ext_clk),
	.D(n2293), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_7__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_7__3_),
	.CK(ext_clk),
	.D(n2292), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_7__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_7__2_),
	.CK(ext_clk),
	.D(n2291), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_7__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_7__1_),
	.CK(ext_clk),
	.D(n2290), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_5__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_5__0_),
	.CK(ext_clk),
	.D(n2281), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_5__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_5__7_),
	.CK(ext_clk),
	.D(n2280), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_5__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_5__6_),
	.CK(ext_clk),
	.D(n2279), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_5__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_5__5_),
	.CK(ext_clk),
	.D(n2278), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_5__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_5__4_),
	.CK(ext_clk),
	.D(n2277), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_5__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_5__2_),
	.CK(ext_clk),
	.D(n2275), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_5__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_5__1_),
	.CK(ext_clk),
	.D(n2274), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_3__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_3__0_),
	.CK(ext_clk),
	.D(n2265), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_3__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_3__7_),
	.CK(ext_clk),
	.D(n2264), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_3__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_3__6_),
	.CK(ext_clk),
	.D(n2263), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_3__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_3__5_),
	.CK(ext_clk),
	.D(n2262), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_3__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_3__4_),
	.CK(ext_clk),
	.D(n2261), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_3__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_3__3_),
	.CK(ext_clk),
	.D(n2260), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_3__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_3__2_),
	.CK(ext_clk),
	.D(n2259), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_3__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_3__1_),
	.CK(ext_clk),
	.D(n2258), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_1__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_1__0_),
	.CK(ext_clk),
	.D(n2249), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_1__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_1__7_),
	.CK(ext_clk),
	.D(n2248), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_1__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_1__6_),
	.CK(ext_clk),
	.D(n2247), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_1__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_1__5_),
	.CK(ext_clk),
	.D(n2246), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_1__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_1__3_),
	.CK(ext_clk),
	.D(n2244), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_1__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_1__2_),
	.CK(ext_clk),
	.D(n2243), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_1__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_1__1_),
	.CK(ext_clk),
	.D(n2242), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_6__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_6__0_),
	.CK(ext_clk),
	.D(n2289), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_6__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_6__7_),
	.CK(ext_clk),
	.D(n2288), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_6__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_6__6_),
	.CK(ext_clk),
	.D(n2287), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_6__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_6__5_),
	.CK(ext_clk),
	.D(n2286), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_6__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_6__4_),
	.CK(ext_clk),
	.D(n2285), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_6__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_6__3_),
	.CK(ext_clk),
	.D(n2284), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_6__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_6__2_),
	.CK(ext_clk),
	.D(n2283), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_6__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_6__1_),
	.CK(ext_clk),
	.D(n2282), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_4__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_4__0_),
	.CK(ext_clk),
	.D(n2273), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_4__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_4__7_),
	.CK(ext_clk),
	.D(n2272), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_4__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_4__6_),
	.CK(ext_clk),
	.D(n2271), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_4__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_4__4_),
	.CK(ext_clk),
	.D(n2269), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_4__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_4__3_),
	.CK(ext_clk),
	.D(n2268), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_4__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_4__2_),
	.CK(ext_clk),
	.D(n2267), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_4__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_4__1_),
	.CK(ext_clk),
	.D(n2266), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_2__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_2__0_),
	.CK(ext_clk),
	.D(n2257), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_2__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_2__7_),
	.CK(ext_clk),
	.D(n2256), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_2__6_ (
	.Q(Mfifo_coe_M_ffmem_mem_2__6_),
	.CK(ext_clk),
	.D(n2255), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_2__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_2__5_),
	.CK(ext_clk),
	.D(n2254), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_2__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_2__4_),
	.CK(ext_clk),
	.D(n2253), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_2__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_2__3_),
	.CK(ext_clk),
	.D(n2252), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_2__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_2__2_),
	.CK(ext_clk),
	.D(n2251), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_2__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_2__1_),
	.CK(ext_clk),
	.D(n2250), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_0__0_ (
	.Q(Mfifo_coe_M_ffmem_mem_0__0_),
	.CK(ext_clk),
	.D(n2241), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_0__7_ (
	.Q(Mfifo_coe_M_ffmem_mem_0__7_),
	.CK(ext_clk),
	.D(n2240), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_0__5_ (
	.Q(Mfifo_coe_M_ffmem_mem_0__5_),
	.CK(ext_clk),
	.D(n2238), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_0__4_ (
	.Q(Mfifo_coe_M_ffmem_mem_0__4_),
	.CK(ext_clk),
	.D(n2237), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_0__3_ (
	.Q(Mfifo_coe_M_ffmem_mem_0__3_),
	.CK(ext_clk),
	.D(n2236), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_0__2_ (
	.Q(Mfifo_coe_M_ffmem_mem_0__2_),
	.CK(ext_clk),
	.D(n2235), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_mem_reg_0__1_ (
	.Q(Mfifo_coe_M_ffmem_mem_0__1_),
	.CK(ext_clk),
	.D(n2234), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_15__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_15__0_),
	.CK(ext_clk),
	.D(n2225), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_15__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_15__7_),
	.CK(ext_clk),
	.D(n2224), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_15__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_15__6_),
	.CK(ext_clk),
	.D(n2223), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_15__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_15__5_),
	.CK(ext_clk),
	.D(n2222), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_15__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_15__4_),
	.CK(ext_clk),
	.D(n2221), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_15__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_15__3_),
	.CK(ext_clk),
	.D(n2220), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_15__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_15__2_),
	.CK(ext_clk),
	.D(n2219), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_15__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_15__1_),
	.CK(ext_clk),
	.D(n2218), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_13__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_13__0_),
	.CK(ext_clk),
	.D(n2209), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_13__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_13__6_),
	.CK(ext_clk),
	.D(n2207), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_13__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_13__5_),
	.CK(ext_clk),
	.D(n2206), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_13__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_13__4_),
	.CK(ext_clk),
	.D(n2205), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_13__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_13__3_),
	.CK(ext_clk),
	.D(n2204), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_13__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_13__2_),
	.CK(ext_clk),
	.D(n2203), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_13__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_13__1_),
	.CK(ext_clk),
	.D(n2202), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_11__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_11__0_),
	.CK(ext_clk),
	.D(n2193), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_11__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_11__7_),
	.CK(ext_clk),
	.D(n2192), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_11__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_11__6_),
	.CK(ext_clk),
	.D(n2191), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_11__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_11__5_),
	.CK(ext_clk),
	.D(n2190), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_11__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_11__4_),
	.CK(ext_clk),
	.D(n2189), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_11__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_11__3_),
	.CK(ext_clk),
	.D(n2188), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_11__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_11__2_),
	.CK(ext_clk),
	.D(n2187), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_11__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_11__1_),
	.CK(ext_clk),
	.D(n2186), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_9__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_9__7_),
	.CK(ext_clk),
	.D(n2176), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_9__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_9__6_),
	.CK(ext_clk),
	.D(n2175), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_9__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_9__5_),
	.CK(ext_clk),
	.D(n2174), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_9__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_9__4_),
	.CK(ext_clk),
	.D(n2173), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_9__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_9__3_),
	.CK(ext_clk),
	.D(n2172), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_9__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_9__2_),
	.CK(ext_clk),
	.D(n2171), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_9__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_9__1_),
	.CK(ext_clk),
	.D(n2170), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_14__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_14__0_),
	.CK(ext_clk),
	.D(n2217), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_14__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_14__7_),
	.CK(ext_clk),
	.D(n2216), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_14__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_14__6_),
	.CK(ext_clk),
	.D(n2215), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_14__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_14__5_),
	.CK(ext_clk),
	.D(n2214), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_14__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_14__4_),
	.CK(ext_clk),
	.D(n2213), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_14__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_14__3_),
	.CK(ext_clk),
	.D(n2212), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_14__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_14__2_),
	.CK(ext_clk),
	.D(n2211), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_12__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_12__0_),
	.CK(ext_clk),
	.D(n2201), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_12__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_12__7_),
	.CK(ext_clk),
	.D(n2200), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_12__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_12__6_),
	.CK(ext_clk),
	.D(n2199), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_12__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_12__5_),
	.CK(ext_clk),
	.D(n2198), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_12__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_12__4_),
	.CK(ext_clk),
	.D(n2197), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_12__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_12__3_),
	.CK(ext_clk),
	.D(n2196), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_12__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_12__2_),
	.CK(ext_clk),
	.D(n2195), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_12__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_12__1_),
	.CK(ext_clk),
	.D(n2194), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_10__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_10__0_),
	.CK(ext_clk),
	.D(n2185), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_10__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_10__7_),
	.CK(ext_clk),
	.D(n2184), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_10__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_10__6_),
	.CK(ext_clk),
	.D(n2183), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_10__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_10__5_),
	.CK(ext_clk),
	.D(n2182), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_10__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_10__4_),
	.CK(ext_clk),
	.D(n2181), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_10__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_10__3_),
	.CK(ext_clk),
	.D(n2180), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_10__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_10__1_),
	.CK(ext_clk),
	.D(n2178), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_8__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_8__0_),
	.CK(ext_clk),
	.D(n2169), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_8__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_8__7_),
	.CK(ext_clk),
	.D(n2168), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_8__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_8__6_),
	.CK(ext_clk),
	.D(n2167), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_8__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_8__5_),
	.CK(ext_clk),
	.D(n2166), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_8__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_8__4_),
	.CK(ext_clk),
	.D(n2165), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_8__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_8__3_),
	.CK(ext_clk),
	.D(n2164), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_8__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_8__2_),
	.CK(ext_clk),
	.D(n2163), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_8__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_8__1_),
	.CK(ext_clk),
	.D(n2162), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_7__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_7__0_),
	.CK(ext_clk),
	.D(n2161), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_7__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_7__7_),
	.CK(ext_clk),
	.D(n2160), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_7__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_7__6_),
	.CK(ext_clk),
	.D(n2159), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_7__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_7__5_),
	.CK(ext_clk),
	.D(n2158), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_7__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_7__4_),
	.CK(ext_clk),
	.D(n2157), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_7__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_7__2_),
	.CK(ext_clk),
	.D(n2155), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_7__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_7__1_),
	.CK(ext_clk),
	.D(n2154), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_5__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_5__0_),
	.CK(ext_clk),
	.D(n2145), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_5__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_5__7_),
	.CK(ext_clk),
	.D(n2144), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_5__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_5__6_),
	.CK(ext_clk),
	.D(n2143), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_5__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_5__5_),
	.CK(ext_clk),
	.D(n2142), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_5__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_5__4_),
	.CK(ext_clk),
	.D(n2141), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_5__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_5__3_),
	.CK(ext_clk),
	.D(n2140), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_5__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_5__2_),
	.CK(ext_clk),
	.D(n2139), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_5__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_5__1_),
	.CK(ext_clk),
	.D(n2138), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_3__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_3__0_),
	.CK(ext_clk),
	.D(n2129), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_3__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_3__7_),
	.CK(ext_clk),
	.D(n2128), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_3__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_3__6_),
	.CK(ext_clk),
	.D(n2127), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_3__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_3__5_),
	.CK(ext_clk),
	.D(n2126), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_3__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_3__3_),
	.CK(ext_clk),
	.D(n2124), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_3__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_3__2_),
	.CK(ext_clk),
	.D(n2123), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_3__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_3__1_),
	.CK(ext_clk),
	.D(n2122), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_1__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_1__0_),
	.CK(ext_clk),
	.D(n2113), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_1__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_1__7_),
	.CK(ext_clk),
	.D(n2112), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_1__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_1__6_),
	.CK(ext_clk),
	.D(n2111), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_1__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_1__5_),
	.CK(ext_clk),
	.D(n2110), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_1__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_1__4_),
	.CK(ext_clk),
	.D(n2109), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_1__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_1__3_),
	.CK(ext_clk),
	.D(n2108), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_1__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_1__2_),
	.CK(ext_clk),
	.D(n2107), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_1__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_1__1_),
	.CK(ext_clk),
	.D(n2106), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_6__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_6__0_),
	.CK(ext_clk),
	.D(n2153), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_6__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_6__7_),
	.CK(ext_clk),
	.D(n2152), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_6__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_6__6_),
	.CK(ext_clk),
	.D(n2151), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_6__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_6__4_),
	.CK(ext_clk),
	.D(n2149), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_6__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_6__3_),
	.CK(ext_clk),
	.D(n2148), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_6__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_6__2_),
	.CK(ext_clk),
	.D(n2147), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_6__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_6__1_),
	.CK(ext_clk),
	.D(n2146), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_4__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_4__0_),
	.CK(ext_clk),
	.D(n2137), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_4__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_4__7_),
	.CK(ext_clk),
	.D(n2136), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_4__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_4__6_),
	.CK(ext_clk),
	.D(n2135), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_4__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_4__5_),
	.CK(ext_clk),
	.D(n2134), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_4__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_4__4_),
	.CK(ext_clk),
	.D(n2133), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_4__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_4__3_),
	.CK(ext_clk),
	.D(n2132), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_4__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_4__2_),
	.CK(ext_clk),
	.D(n2131), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_4__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_4__1_),
	.CK(ext_clk),
	.D(n2130), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_2__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_2__0_),
	.CK(ext_clk),
	.D(n2121), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_2__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_2__7_),
	.CK(ext_clk),
	.D(n2120), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_2__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_2__5_),
	.CK(ext_clk),
	.D(n2118), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_2__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_2__4_),
	.CK(ext_clk),
	.D(n2117), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_2__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_2__3_),
	.CK(ext_clk),
	.D(n2116), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_2__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_2__2_),
	.CK(ext_clk),
	.D(n2115), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_2__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_2__1_),
	.CK(ext_clk),
	.D(n2114), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_0__0_ (
	.Q(Mfifo_xin_M_ffmem_mem_0__0_),
	.CK(ext_clk),
	.D(n2105), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_0__7_ (
	.Q(Mfifo_xin_M_ffmem_mem_0__7_),
	.CK(ext_clk),
	.D(n2104), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_0__6_ (
	.Q(Mfifo_xin_M_ffmem_mem_0__6_),
	.CK(ext_clk),
	.D(n2103), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_0__5_ (
	.Q(Mfifo_xin_M_ffmem_mem_0__5_),
	.CK(ext_clk),
	.D(n2102), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_0__4_ (
	.Q(Mfifo_xin_M_ffmem_mem_0__4_),
	.CK(ext_clk),
	.D(n2101), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_0__3_ (
	.Q(Mfifo_xin_M_ffmem_mem_0__3_),
	.CK(ext_clk),
	.D(n2100), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_0__2_ (
	.Q(Mfifo_xin_M_ffmem_mem_0__2_),
	.CK(ext_clk),
	.D(n2099), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_mem_reg_0__1_ (
	.Q(Mfifo_xin_M_ffmem_mem_0__1_),
	.CK(ext_clk),
	.D(n2098), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_rdata_reg_2_ (
	.Q(int_coe[2]),
	.CK(int_clk),
	.D(n2232), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_rdata_reg_5_ (
	.Q(int_coe[5]),
	.CK(int_clk),
	.D(n2229), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_coe_M_ffmem_rdata_reg_6_ (
	.Q(int_coe[6]),
	.CK(int_clk),
	.D(n2228), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_rdata_reg_1_ (
	.Q(int_xin[1]),
	.CK(int_clk),
	.D(n2097), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_rdata_reg_2_ (
	.Q(int_xin[2]),
	.CK(int_clk),
	.D(n2096), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_rdata_reg_3_ (
	.Q(int_xin[3]),
	.CK(int_clk),
	.D(n2095), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_rdata_reg_4_ (
	.Q(int_xin[4]),
	.CK(int_clk),
	.D(n2094), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_rdata_reg_5_ (
	.Q(int_xin[5]),
	.CK(int_clk),
	.D(n2093), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_rdata_reg_6_ (
	.Q(int_xin[6]),
	.CK(int_clk),
	.D(n2092), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_rdata_reg_7_ (
	.Q(int_xin[7]),
	.CK(int_clk),
	.D(n2091), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_xin_M_ffmem_rdata_reg_0_ (
	.Q(int_xin[0]),
	.CK(int_clk),
	.D(n2090), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__21_),
	.CK(int_clk),
	.D(n2064), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__21_),
	.CK(int_clk),
	.D(n2063), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__21_),
	.CK(int_clk),
	.D(n2062), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__21_),
	.CK(int_clk),
	.D(n2061), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__21_),
	.CK(int_clk),
	.D(n2060), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__21_),
	.CK(int_clk),
	.D(n2059), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__21_),
	.CK(int_clk),
	.D(n2058), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__21_),
	.CK(int_clk),
	.D(n2057), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__21_),
	.CK(int_clk),
	.D(n2056), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__21_),
	.CK(int_clk),
	.D(n2055), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__21_),
	.CK(int_clk),
	.D(n2054), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__21_),
	.CK(int_clk),
	.D(n2053), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__21_),
	.CK(int_clk),
	.D(n2052), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__21_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__21_),
	.CK(int_clk),
	.D(n2051), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__22_),
	.CK(int_clk),
	.D(n2049), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__22_),
	.CK(int_clk),
	.D(n2048), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__22_),
	.CK(int_clk),
	.D(n2047), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__22_),
	.CK(int_clk),
	.D(n2046), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__22_),
	.CK(int_clk),
	.D(n2045), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__22_),
	.CK(int_clk),
	.D(n2044), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__22_),
	.CK(int_clk),
	.D(n2043), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__22_),
	.CK(int_clk),
	.D(n2042), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__22_),
	.CK(int_clk),
	.D(n2041), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__22_),
	.CK(int_clk),
	.D(n2040), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__22_),
	.CK(int_clk),
	.D(n2039), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__22_),
	.CK(int_clk),
	.D(n2038), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__22_),
	.CK(int_clk),
	.D(n2037), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__22_),
	.CK(int_clk),
	.D(n2036), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__22_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__22_),
	.CK(int_clk),
	.D(n2034), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__23_),
	.CK(int_clk),
	.D(n2033), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__23_),
	.CK(int_clk),
	.D(n2032), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__23_),
	.CK(int_clk),
	.D(n2031), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__23_),
	.CK(int_clk),
	.D(n2030), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__23_),
	.CK(int_clk),
	.D(n2029), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__23_),
	.CK(int_clk),
	.D(n2028), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__23_),
	.CK(int_clk),
	.D(n2027), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__23_),
	.CK(int_clk),
	.D(n2026), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__23_),
	.CK(int_clk),
	.D(n2025), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__23_),
	.CK(int_clk),
	.D(n2024), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__23_),
	.CK(int_clk),
	.D(n2023), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__23_),
	.CK(int_clk),
	.D(n2022), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__23_),
	.CK(int_clk),
	.D(n2021), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__23_),
	.CK(int_clk),
	.D(n2019), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__23_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__23_),
	.CK(int_clk),
	.D(n2018), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__24_),
	.CK(int_clk),
	.D(n2017), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__24_),
	.CK(int_clk),
	.D(n2016), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__24_),
	.CK(int_clk),
	.D(n2015), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__24_),
	.CK(int_clk),
	.D(n2014), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__24_),
	.CK(int_clk),
	.D(n2013), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__24_),
	.CK(int_clk),
	.D(n2012), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__24_),
	.CK(int_clk),
	.D(n2011), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__24_),
	.CK(int_clk),
	.D(n2010), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__24_),
	.CK(int_clk),
	.D(n2009), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__24_),
	.CK(int_clk),
	.D(n2008), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__24_),
	.CK(int_clk),
	.D(n2007), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__24_),
	.CK(int_clk),
	.D(n2006), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__24_),
	.CK(int_clk),
	.D(n2004), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__24_),
	.CK(int_clk),
	.D(n2003), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__24_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__24_),
	.CK(int_clk),
	.D(n2002), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__25_),
	.CK(int_clk),
	.D(n2001), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__25_),
	.CK(int_clk),
	.D(n2000), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__25_),
	.CK(int_clk),
	.D(n1999), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__25_),
	.CK(int_clk),
	.D(n1998), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__25_),
	.CK(int_clk),
	.D(n1997), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__25_),
	.CK(int_clk),
	.D(n1996), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__25_),
	.CK(int_clk),
	.D(n1995), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__25_),
	.CK(int_clk),
	.D(n1994), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__25_),
	.CK(int_clk),
	.D(n1993), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__25_),
	.CK(int_clk),
	.D(n1992), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__25_),
	.CK(int_clk),
	.D(n1991), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__25_),
	.CK(int_clk),
	.D(n1989), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__25_),
	.CK(int_clk),
	.D(n1988), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__25_),
	.CK(int_clk),
	.D(n1987), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__25_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__25_),
	.CK(int_clk),
	.D(n1986), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__26_),
	.CK(int_clk),
	.D(n1985), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__26_),
	.CK(int_clk),
	.D(n1984), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__26_),
	.CK(int_clk),
	.D(n1983), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__26_),
	.CK(int_clk),
	.D(n1982), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__26_),
	.CK(int_clk),
	.D(n1981), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__26_),
	.CK(int_clk),
	.D(n1980), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__26_),
	.CK(int_clk),
	.D(n1979), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__26_),
	.CK(int_clk),
	.D(n1978), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__26_),
	.CK(int_clk),
	.D(n1977), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__26_),
	.CK(int_clk),
	.D(n1976), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__26_),
	.CK(int_clk),
	.D(n1974), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__26_),
	.CK(int_clk),
	.D(n1973), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__26_),
	.CK(int_clk),
	.D(n1972), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__26_),
	.CK(int_clk),
	.D(n1971), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__26_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__26_),
	.CK(int_clk),
	.D(n1970), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__27_),
	.CK(int_clk),
	.D(n1969), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__27_),
	.CK(int_clk),
	.D(n1968), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__27_),
	.CK(int_clk),
	.D(n1967), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__27_),
	.CK(int_clk),
	.D(n1966), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__27_),
	.CK(int_clk),
	.D(n1965), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__27_),
	.CK(int_clk),
	.D(n1964), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__27_),
	.CK(int_clk),
	.D(n1963), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__27_),
	.CK(int_clk),
	.D(n1962), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__27_),
	.CK(int_clk),
	.D(n1961), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__27_),
	.CK(int_clk),
	.D(n1959), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__27_),
	.CK(int_clk),
	.D(n1958), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__27_),
	.CK(int_clk),
	.D(n1957), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__27_),
	.CK(int_clk),
	.D(n1956), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__27_),
	.CK(int_clk),
	.D(n1955), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__27_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__27_),
	.CK(int_clk),
	.D(n1954), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__28_),
	.CK(int_clk),
	.D(n1953), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__28_),
	.CK(int_clk),
	.D(n1952), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__28_),
	.CK(int_clk),
	.D(n1951), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__28_),
	.CK(int_clk),
	.D(n1950), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__28_),
	.CK(int_clk),
	.D(n1949), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__28_),
	.CK(int_clk),
	.D(n1948), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__28_),
	.CK(int_clk),
	.D(n1947), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__28_),
	.CK(int_clk),
	.D(n1946), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__28_),
	.CK(int_clk),
	.D(n1944), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__28_),
	.CK(int_clk),
	.D(n1943), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__28_),
	.CK(int_clk),
	.D(n1942), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__28_),
	.CK(int_clk),
	.D(n1941), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__28_),
	.CK(int_clk),
	.D(n1940), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__28_),
	.CK(int_clk),
	.D(n1939), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__28_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__28_),
	.CK(int_clk),
	.D(n1938), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__29_),
	.CK(int_clk),
	.D(n1937), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__29_),
	.CK(int_clk),
	.D(n1936), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__29_),
	.CK(int_clk),
	.D(n1935), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__29_),
	.CK(int_clk),
	.D(n1934), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__29_),
	.CK(int_clk),
	.D(n1933), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__29_),
	.CK(int_clk),
	.D(n1932), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__29_),
	.CK(int_clk),
	.D(n1931), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__29_),
	.CK(int_clk),
	.D(n1929), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__29_),
	.CK(int_clk),
	.D(n1928), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__29_),
	.CK(int_clk),
	.D(n1927), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__29_),
	.CK(int_clk),
	.D(n1926), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__29_),
	.CK(int_clk),
	.D(n1925), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__29_),
	.CK(int_clk),
	.D(n1924), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__29_),
	.CK(int_clk),
	.D(n1923), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__29_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__29_),
	.CK(int_clk),
	.D(n1922), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__30_),
	.CK(int_clk),
	.D(n1921), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__30_),
	.CK(int_clk),
	.D(n1920), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__30_),
	.CK(int_clk),
	.D(n1919), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__30_),
	.CK(int_clk),
	.D(n1918), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__30_),
	.CK(int_clk),
	.D(n1917), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__30_),
	.CK(int_clk),
	.D(n1916), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__30_),
	.CK(int_clk),
	.D(n1914), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__30_),
	.CK(int_clk),
	.D(n1913), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__30_),
	.CK(int_clk),
	.D(n1912), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__30_),
	.CK(int_clk),
	.D(n1911), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__30_),
	.CK(int_clk),
	.D(n1910), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__30_),
	.CK(int_clk),
	.D(n1909), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__30_),
	.CK(int_clk),
	.D(n1908), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__30_),
	.CK(int_clk),
	.D(n1907), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__30_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__30_),
	.CK(int_clk),
	.D(n1906), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__31_),
	.CK(int_clk),
	.D(n1905), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__31_),
	.CK(int_clk),
	.D(n1904), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__31_),
	.CK(int_clk),
	.D(n1903), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__31_),
	.CK(int_clk),
	.D(n1902), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__31_),
	.CK(int_clk),
	.D(n1901), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__31_),
	.CK(int_clk),
	.D(n1899), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__31_),
	.CK(int_clk),
	.D(n1898), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__31_),
	.CK(int_clk),
	.D(n1897), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__31_),
	.CK(int_clk),
	.D(n1896), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__31_),
	.CK(int_clk),
	.D(n1895), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__31_),
	.CK(int_clk),
	.D(n1894), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__31_),
	.CK(int_clk),
	.D(n1893), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__31_),
	.CK(int_clk),
	.D(n1892), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__31_),
	.CK(int_clk),
	.D(n1891), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__31_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__31_),
	.CK(int_clk),
	.D(n1890), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__32_),
	.CK(int_clk),
	.D(n1889), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__32_),
	.CK(int_clk),
	.D(n1888), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__32_),
	.CK(int_clk),
	.D(n1887), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__32_),
	.CK(int_clk),
	.D(n1886), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__32_),
	.CK(int_clk),
	.D(n1884), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__32_),
	.CK(int_clk),
	.D(n1883), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__32_),
	.CK(int_clk),
	.D(n1882), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__32_),
	.CK(int_clk),
	.D(n1881), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__32_),
	.CK(int_clk),
	.D(n1880), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__32_),
	.CK(int_clk),
	.D(n1879), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__32_),
	.CK(int_clk),
	.D(n1878), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__32_),
	.CK(int_clk),
	.D(n1877), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__32_),
	.CK(int_clk),
	.D(n1876), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__32_),
	.CK(int_clk),
	.D(n1875), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__32_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__32_),
	.CK(int_clk),
	.D(n1874), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__33_),
	.CK(int_clk),
	.D(n1873), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__33_),
	.CK(int_clk),
	.D(n1872), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__33_),
	.CK(int_clk),
	.D(n1871), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__33_),
	.CK(int_clk),
	.D(n1869), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__33_),
	.CK(int_clk),
	.D(n1868), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__33_),
	.CK(int_clk),
	.D(n1867), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__33_),
	.CK(int_clk),
	.D(n1866), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__33_),
	.CK(int_clk),
	.D(n1865), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__33_),
	.CK(int_clk),
	.D(n1864), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__33_),
	.CK(int_clk),
	.D(n1863), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__33_),
	.CK(int_clk),
	.D(n1862), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__33_),
	.CK(int_clk),
	.D(n1861), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__33_),
	.CK(int_clk),
	.D(n1860), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__33_),
	.CK(int_clk),
	.D(n1859), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__33_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__33_),
	.CK(int_clk),
	.D(n1858), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__34_),
	.CK(int_clk),
	.D(n1857), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__34_),
	.CK(int_clk),
	.D(n1856), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__34_),
	.CK(int_clk),
	.D(n1854), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__34_),
	.CK(int_clk),
	.D(n1853), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__34_),
	.CK(int_clk),
	.D(n1852), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__34_),
	.CK(int_clk),
	.D(n1851), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__34_),
	.CK(int_clk),
	.D(n1850), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__34_),
	.CK(int_clk),
	.D(n1849), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__34_),
	.CK(int_clk),
	.D(n1848), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__34_),
	.CK(int_clk),
	.D(n1847), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__34_),
	.CK(int_clk),
	.D(n1846), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__34_),
	.CK(int_clk),
	.D(n1845), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__34_),
	.CK(int_clk),
	.D(n1844), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__34_),
	.CK(int_clk),
	.D(n1843), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__34_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__34_),
	.CK(int_clk),
	.D(n1842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__35_),
	.CK(int_clk),
	.D(n1841), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__35_),
	.CK(int_clk),
	.D(n1839), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__35_),
	.CK(int_clk),
	.D(n1838), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__35_),
	.CK(int_clk),
	.D(n1837), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__35_),
	.CK(int_clk),
	.D(n1836), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__35_),
	.CK(int_clk),
	.D(n1835), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__35_),
	.CK(int_clk),
	.D(n1834), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__35_),
	.CK(int_clk),
	.D(n1833), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__35_),
	.CK(int_clk),
	.D(n1832), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__35_),
	.CK(int_clk),
	.D(n1831), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__35_),
	.CK(int_clk),
	.D(n1830), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__35_),
	.CK(int_clk),
	.D(n1829), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__35_),
	.CK(int_clk),
	.D(n1828), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__35_),
	.CK(int_clk),
	.D(n1827), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__35_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__35_),
	.CK(int_clk),
	.D(n1826), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__36_),
	.CK(int_clk),
	.D(n1824), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__36_),
	.CK(int_clk),
	.D(n1823), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__36_),
	.CK(int_clk),
	.D(n1822), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__36_),
	.CK(int_clk),
	.D(n1821), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__36_),
	.CK(int_clk),
	.D(n1820), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__36_),
	.CK(int_clk),
	.D(n1819), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__36_),
	.CK(int_clk),
	.D(n1818), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__36_),
	.CK(int_clk),
	.D(n1817), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__36_),
	.CK(int_clk),
	.D(n1816), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__36_),
	.CK(int_clk),
	.D(n1815), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__36_),
	.CK(int_clk),
	.D(n1814), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__36_),
	.CK(int_clk),
	.D(n1813), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__36_),
	.CK(int_clk),
	.D(n1812), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__36_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__36_),
	.CK(int_clk),
	.D(n1811), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__37_),
	.CK(int_clk),
	.D(n1809), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__37_),
	.CK(int_clk),
	.D(n1808), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__37_),
	.CK(int_clk),
	.D(n1807), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__37_),
	.CK(int_clk),
	.D(n1806), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__37_),
	.CK(int_clk),
	.D(n1805), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__37_),
	.CK(int_clk),
	.D(n1804), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__37_),
	.CK(int_clk),
	.D(n1803), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__37_),
	.CK(int_clk),
	.D(n1802), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__37_),
	.CK(int_clk),
	.D(n1801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__37_),
	.CK(int_clk),
	.D(n1800), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__37_),
	.CK(int_clk),
	.D(n1799), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__37_),
	.CK(int_clk),
	.D(n1798), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__37_),
	.CK(int_clk),
	.D(n1797), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__37_),
	.CK(int_clk),
	.D(n1796), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__37_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__37_),
	.CK(int_clk),
	.D(n1794), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__38_),
	.CK(int_clk),
	.D(n1793), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__38_),
	.CK(int_clk),
	.D(n1792), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__38_),
	.CK(int_clk),
	.D(n1791), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__38_),
	.CK(int_clk),
	.D(n1790), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__38_),
	.CK(int_clk),
	.D(n1789), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__38_),
	.CK(int_clk),
	.D(n1788), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__38_),
	.CK(int_clk),
	.D(n1787), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__38_),
	.CK(int_clk),
	.D(n1786), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__38_),
	.CK(int_clk),
	.D(n1785), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__38_),
	.CK(int_clk),
	.D(n1784), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__38_),
	.CK(int_clk),
	.D(n1783), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__38_),
	.CK(int_clk),
	.D(n1782), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__38_),
	.CK(int_clk),
	.D(n1781), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__38_),
	.CK(int_clk),
	.D(n1779), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__38_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__38_),
	.CK(int_clk),
	.D(n1778), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__39_),
	.CK(int_clk),
	.D(n1777), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__39_),
	.CK(int_clk),
	.D(n1776), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__39_),
	.CK(int_clk),
	.D(n1775), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__39_),
	.CK(int_clk),
	.D(n1774), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__39_),
	.CK(int_clk),
	.D(n1773), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__39_),
	.CK(int_clk),
	.D(n1772), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__39_),
	.CK(int_clk),
	.D(n1771), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__39_),
	.CK(int_clk),
	.D(n1770), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__39_),
	.CK(int_clk),
	.D(n1769), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__39_),
	.CK(int_clk),
	.D(n1768), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__39_),
	.CK(int_clk),
	.D(n1767), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__39_),
	.CK(int_clk),
	.D(n1766), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__39_),
	.CK(int_clk),
	.D(n1764), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__39_),
	.CK(int_clk),
	.D(n1763), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__39_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__39_),
	.CK(int_clk),
	.D(n1762), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__40_),
	.CK(int_clk),
	.D(n1761), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__40_),
	.CK(int_clk),
	.D(n1760), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__40_),
	.CK(int_clk),
	.D(n1759), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__40_),
	.CK(int_clk),
	.D(n1758), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__40_),
	.CK(int_clk),
	.D(n1757), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__40_),
	.CK(int_clk),
	.D(n1756), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__40_),
	.CK(int_clk),
	.D(n1755), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__40_),
	.CK(int_clk),
	.D(n1754), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__40_),
	.CK(int_clk),
	.D(n1753), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__40_),
	.CK(int_clk),
	.D(n1752), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__40_),
	.CK(int_clk),
	.D(n1751), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__40_),
	.CK(int_clk),
	.D(n1749), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__40_),
	.CK(int_clk),
	.D(n1748), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__40_),
	.CK(int_clk),
	.D(n1747), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__40_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__40_),
	.CK(int_clk),
	.D(n1746), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__41_),
	.CK(int_clk),
	.D(n1745), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__41_),
	.CK(int_clk),
	.D(n1744), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__41_),
	.CK(int_clk),
	.D(n1743), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__41_),
	.CK(int_clk),
	.D(n1742), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__41_),
	.CK(int_clk),
	.D(n1741), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__41_),
	.CK(int_clk),
	.D(n1740), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__41_),
	.CK(int_clk),
	.D(n1739), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__41_),
	.CK(int_clk),
	.D(n1738), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__41_),
	.CK(int_clk),
	.D(n1737), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__41_),
	.CK(int_clk),
	.D(n1736), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__41_),
	.CK(int_clk),
	.D(n1734), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__41_),
	.CK(int_clk),
	.D(n1733), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__41_),
	.CK(int_clk),
	.D(n1732), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__41_),
	.CK(int_clk),
	.D(n1731), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__41_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__41_),
	.CK(int_clk),
	.D(n1730), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__0_),
	.CK(int_clk),
	.D(n1729), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__0_),
	.CK(int_clk),
	.D(n1728), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__0_),
	.CK(int_clk),
	.D(n1727), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__0_),
	.CK(int_clk),
	.D(n1726), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__0_),
	.CK(int_clk),
	.D(n1725), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__0_),
	.CK(int_clk),
	.D(n1724), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__0_),
	.CK(int_clk),
	.D(n1723), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__0_),
	.CK(int_clk),
	.D(n1722), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__0_),
	.CK(int_clk),
	.D(n1721), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__0_),
	.CK(int_clk),
	.D(n1719), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__0_),
	.CK(int_clk),
	.D(n1718), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__0_),
	.CK(int_clk),
	.D(n1717), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__0_),
	.CK(int_clk),
	.D(n1716), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__0_),
	.CK(int_clk),
	.D(n1715), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__0_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__0_),
	.CK(int_clk),
	.D(n1714), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__1_),
	.CK(int_clk),
	.D(n1713), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__1_),
	.CK(int_clk),
	.D(n1712), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__1_),
	.CK(int_clk),
	.D(n1711), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__1_),
	.CK(int_clk),
	.D(n1710), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__1_),
	.CK(int_clk),
	.D(n1709), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__1_),
	.CK(int_clk),
	.D(n1708), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__1_),
	.CK(int_clk),
	.D(n1707), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__1_),
	.CK(int_clk),
	.D(n1706), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__1_),
	.CK(int_clk),
	.D(n1704), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__1_),
	.CK(int_clk),
	.D(n1703), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__1_),
	.CK(int_clk),
	.D(n1702), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__1_),
	.CK(int_clk),
	.D(n1701), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__1_),
	.CK(int_clk),
	.D(n1700), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__1_),
	.CK(int_clk),
	.D(n1699), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__1_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__1_),
	.CK(int_clk),
	.D(n1698), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__2_),
	.CK(int_clk),
	.D(n1697), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__2_),
	.CK(int_clk),
	.D(n1696), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__2_),
	.CK(int_clk),
	.D(n1695), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__2_),
	.CK(int_clk),
	.D(n1694), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__2_),
	.CK(int_clk),
	.D(n1693), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__2_),
	.CK(int_clk),
	.D(n1692), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__2_),
	.CK(int_clk),
	.D(n1691), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__2_),
	.CK(int_clk),
	.D(n1689), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__2_),
	.CK(int_clk),
	.D(n1688), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__2_),
	.CK(int_clk),
	.D(n1687), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__2_),
	.CK(int_clk),
	.D(n1686), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__2_),
	.CK(int_clk),
	.D(n1685), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__2_),
	.CK(int_clk),
	.D(n1684), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__2_),
	.CK(int_clk),
	.D(n1683), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__2_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__2_),
	.CK(int_clk),
	.D(n1682), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__3_),
	.CK(int_clk),
	.D(n1681), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__3_),
	.CK(int_clk),
	.D(n1680), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__3_),
	.CK(int_clk),
	.D(n1679), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__3_),
	.CK(int_clk),
	.D(n1678), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__3_),
	.CK(int_clk),
	.D(n1677), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__3_),
	.CK(int_clk),
	.D(n1676), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__3_),
	.CK(int_clk),
	.D(n1674), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__3_),
	.CK(int_clk),
	.D(n1673), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__3_),
	.CK(int_clk),
	.D(n1672), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__3_),
	.CK(int_clk),
	.D(n1671), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__3_),
	.CK(int_clk),
	.D(n1670), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__3_),
	.CK(int_clk),
	.D(n1669), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__3_),
	.CK(int_clk),
	.D(n1668), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__3_),
	.CK(int_clk),
	.D(n1667), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__3_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__3_),
	.CK(int_clk),
	.D(n1666), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__4_),
	.CK(int_clk),
	.D(n1665), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__4_),
	.CK(int_clk),
	.D(n1664), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__4_),
	.CK(int_clk),
	.D(n1663), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__4_),
	.CK(int_clk),
	.D(n1662), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__4_),
	.CK(int_clk),
	.D(n1661), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__4_),
	.CK(int_clk),
	.D(n1659), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__4_),
	.CK(int_clk),
	.D(n1658), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__4_),
	.CK(int_clk),
	.D(n1657), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__4_),
	.CK(int_clk),
	.D(n1656), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__4_),
	.CK(int_clk),
	.D(n1655), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__4_),
	.CK(int_clk),
	.D(n1654), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__4_),
	.CK(int_clk),
	.D(n1653), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__4_),
	.CK(int_clk),
	.D(n1652), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__4_),
	.CK(int_clk),
	.D(n1651), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__4_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__4_),
	.CK(int_clk),
	.D(n1650), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__5_),
	.CK(int_clk),
	.D(n1649), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__5_),
	.CK(int_clk),
	.D(n1648), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__5_),
	.CK(int_clk),
	.D(n1647), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__5_),
	.CK(int_clk),
	.D(n1646), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__5_),
	.CK(int_clk),
	.D(n1644), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__5_),
	.CK(int_clk),
	.D(n1643), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__5_),
	.CK(int_clk),
	.D(n1642), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__5_),
	.CK(int_clk),
	.D(n1641), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__5_),
	.CK(int_clk),
	.D(n1640), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__5_),
	.CK(int_clk),
	.D(n1639), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__5_),
	.CK(int_clk),
	.D(n1638), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__5_),
	.CK(int_clk),
	.D(n1637), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__5_),
	.CK(int_clk),
	.D(n1636), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__5_),
	.CK(int_clk),
	.D(n1635), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__5_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__5_),
	.CK(int_clk),
	.D(n1634), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__6_),
	.CK(int_clk),
	.D(n1633), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__6_),
	.CK(int_clk),
	.D(n1632), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__6_),
	.CK(int_clk),
	.D(n1631), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__6_),
	.CK(int_clk),
	.D(n1629), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__6_),
	.CK(int_clk),
	.D(n1628), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__6_),
	.CK(int_clk),
	.D(n1627), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__6_),
	.CK(int_clk),
	.D(n1626), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__6_),
	.CK(int_clk),
	.D(n1625), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__6_),
	.CK(int_clk),
	.D(n1624), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__6_),
	.CK(int_clk),
	.D(n1623), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__6_),
	.CK(int_clk),
	.D(n1622), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__6_),
	.CK(int_clk),
	.D(n1621), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__6_),
	.CK(int_clk),
	.D(n1620), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__6_),
	.CK(int_clk),
	.D(n1619), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__6_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__6_),
	.CK(int_clk),
	.D(n1618), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__7_),
	.CK(int_clk),
	.D(n1617), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__7_),
	.CK(int_clk),
	.D(n1616), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__7_),
	.CK(int_clk),
	.D(n1614), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__7_),
	.CK(int_clk),
	.D(n1613), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__7_),
	.CK(int_clk),
	.D(n1612), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__7_),
	.CK(int_clk),
	.D(n1611), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__7_),
	.CK(int_clk),
	.D(n1610), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__7_),
	.CK(int_clk),
	.D(n1609), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__7_),
	.CK(int_clk),
	.D(n1608), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__7_),
	.CK(int_clk),
	.D(n1607), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__7_),
	.CK(int_clk),
	.D(n1606), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__7_),
	.CK(int_clk),
	.D(n1605), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__7_),
	.CK(int_clk),
	.D(n1604), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__7_),
	.CK(int_clk),
	.D(n1603), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__7_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__7_),
	.CK(int_clk),
	.D(n1602), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__8_),
	.CK(int_clk),
	.D(n1601), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__8_),
	.CK(int_clk),
	.D(n1599), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__8_),
	.CK(int_clk),
	.D(n1598), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__8_),
	.CK(int_clk),
	.D(n1597), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__8_),
	.CK(int_clk),
	.D(n1596), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__8_),
	.CK(int_clk),
	.D(n1595), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__8_),
	.CK(int_clk),
	.D(n1594), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__8_),
	.CK(int_clk),
	.D(n1593), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__8_),
	.CK(int_clk),
	.D(n1592), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__8_),
	.CK(int_clk),
	.D(n1591), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__8_),
	.CK(int_clk),
	.D(n1590), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__8_),
	.CK(int_clk),
	.D(n1589), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__8_),
	.CK(int_clk),
	.D(n1588), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__8_),
	.CK(int_clk),
	.D(n1587), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__8_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__8_),
	.CK(int_clk),
	.D(n1586), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__9_),
	.CK(int_clk),
	.D(n1584), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__9_),
	.CK(int_clk),
	.D(n1583), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__9_),
	.CK(int_clk),
	.D(n1582), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__9_),
	.CK(int_clk),
	.D(n1581), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__9_),
	.CK(int_clk),
	.D(n1580), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__9_),
	.CK(int_clk),
	.D(n1579), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__9_),
	.CK(int_clk),
	.D(n1578), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__9_),
	.CK(int_clk),
	.D(n1577), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__9_),
	.CK(int_clk),
	.D(n1576), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__9_),
	.CK(int_clk),
	.D(n1575), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__9_),
	.CK(int_clk),
	.D(n1574), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__9_),
	.CK(int_clk),
	.D(n1573), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__9_),
	.CK(int_clk),
	.D(n1572), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__9_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__9_),
	.CK(int_clk),
	.D(n1571), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__10_),
	.CK(int_clk),
	.D(n1569), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__10_),
	.CK(int_clk),
	.D(n1568), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__10_),
	.CK(int_clk),
	.D(n1567), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__10_),
	.CK(int_clk),
	.D(n1566), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__10_),
	.CK(int_clk),
	.D(n1565), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__10_),
	.CK(int_clk),
	.D(n1564), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__10_),
	.CK(int_clk),
	.D(n1563), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__10_),
	.CK(int_clk),
	.D(n1562), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__10_),
	.CK(int_clk),
	.D(n1561), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__10_),
	.CK(int_clk),
	.D(n1560), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__10_),
	.CK(int_clk),
	.D(n1559), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__10_),
	.CK(int_clk),
	.D(n1558), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__10_),
	.CK(int_clk),
	.D(n1557), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__10_),
	.CK(int_clk),
	.D(n1556), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__10_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__10_),
	.CK(int_clk),
	.D(n1554), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__11_),
	.CK(int_clk),
	.D(n1553), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__11_),
	.CK(int_clk),
	.D(n1552), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__11_),
	.CK(int_clk),
	.D(n1551), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__11_),
	.CK(int_clk),
	.D(n1550), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__11_),
	.CK(int_clk),
	.D(n1549), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__11_),
	.CK(int_clk),
	.D(n1548), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__11_),
	.CK(int_clk),
	.D(n1547), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__11_),
	.CK(int_clk),
	.D(n1546), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__11_),
	.CK(int_clk),
	.D(n1545), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__11_),
	.CK(int_clk),
	.D(n1544), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__11_),
	.CK(int_clk),
	.D(n1543), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__11_),
	.CK(int_clk),
	.D(n1542), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__11_),
	.CK(int_clk),
	.D(n1541), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__11_),
	.CK(int_clk),
	.D(n1539), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__11_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__11_),
	.CK(int_clk),
	.D(n1538), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__12_),
	.CK(int_clk),
	.D(n1537), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__12_),
	.CK(int_clk),
	.D(n1536), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__12_),
	.CK(int_clk),
	.D(n1535), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__12_),
	.CK(int_clk),
	.D(n1534), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__12_),
	.CK(int_clk),
	.D(n1533), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__12_),
	.CK(int_clk),
	.D(n1532), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__12_),
	.CK(int_clk),
	.D(n1531), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__12_),
	.CK(int_clk),
	.D(n1530), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__12_),
	.CK(int_clk),
	.D(n1529), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__12_),
	.CK(int_clk),
	.D(n1528), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__12_),
	.CK(int_clk),
	.D(n1527), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__12_),
	.CK(int_clk),
	.D(n1526), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__12_),
	.CK(int_clk),
	.D(n1524), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__12_),
	.CK(int_clk),
	.D(n1523), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__12_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__12_),
	.CK(int_clk),
	.D(n1522), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__13_),
	.CK(int_clk),
	.D(n1521), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__13_),
	.CK(int_clk),
	.D(n1520), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__13_),
	.CK(int_clk),
	.D(n1519), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__13_),
	.CK(int_clk),
	.D(n1518), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__13_),
	.CK(int_clk),
	.D(n1517), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__13_),
	.CK(int_clk),
	.D(n1516), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__13_),
	.CK(int_clk),
	.D(n1515), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__13_),
	.CK(int_clk),
	.D(n1514), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__13_),
	.CK(int_clk),
	.D(n1513), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__13_),
	.CK(int_clk),
	.D(n1512), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__13_),
	.CK(int_clk),
	.D(n1511), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__13_),
	.CK(int_clk),
	.D(n1509), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__13_),
	.CK(int_clk),
	.D(n1508), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__13_),
	.CK(int_clk),
	.D(n1507), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__13_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__13_),
	.CK(int_clk),
	.D(n1506), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__14_),
	.CK(int_clk),
	.D(n1505), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__14_),
	.CK(int_clk),
	.D(n1504), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__14_),
	.CK(int_clk),
	.D(n1503), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__14_),
	.CK(int_clk),
	.D(n1502), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__14_),
	.CK(int_clk),
	.D(n1501), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__14_),
	.CK(int_clk),
	.D(n1500), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__14_),
	.CK(int_clk),
	.D(n1499), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__14_),
	.CK(int_clk),
	.D(n1498), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__14_),
	.CK(int_clk),
	.D(n1497), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__14_),
	.CK(int_clk),
	.D(n1496), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__14_),
	.CK(int_clk),
	.D(n1494), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__14_),
	.CK(int_clk),
	.D(n1493), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__14_),
	.CK(int_clk),
	.D(n1492), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__14_),
	.CK(int_clk),
	.D(n1491), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__14_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__14_),
	.CK(int_clk),
	.D(n1490), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__15_),
	.CK(int_clk),
	.D(n1489), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__15_),
	.CK(int_clk),
	.D(n1488), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__15_),
	.CK(int_clk),
	.D(n1487), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__15_),
	.CK(int_clk),
	.D(n1486), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__15_),
	.CK(int_clk),
	.D(n1485), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__15_),
	.CK(int_clk),
	.D(n1484), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__15_),
	.CK(int_clk),
	.D(n1483), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__15_),
	.CK(int_clk),
	.D(n1482), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__15_),
	.CK(int_clk),
	.D(n1481), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__15_),
	.CK(int_clk),
	.D(n1479), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__15_),
	.CK(int_clk),
	.D(n1478), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__15_),
	.CK(int_clk),
	.D(n1477), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__15_),
	.CK(int_clk),
	.D(n1476), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__15_),
	.CK(int_clk),
	.D(n1475), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__15_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__15_),
	.CK(int_clk),
	.D(n1474), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__16_),
	.CK(int_clk),
	.D(n1473), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__16_),
	.CK(int_clk),
	.D(n1472), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__16_),
	.CK(int_clk),
	.D(n1471), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__16_),
	.CK(int_clk),
	.D(n1470), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__16_),
	.CK(int_clk),
	.D(n1469), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__16_),
	.CK(int_clk),
	.D(n1468), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__16_),
	.CK(int_clk),
	.D(n1467), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__16_),
	.CK(int_clk),
	.D(n1466), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__16_),
	.CK(int_clk),
	.D(n1464), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__16_),
	.CK(int_clk),
	.D(n1463), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__16_),
	.CK(int_clk),
	.D(n1462), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__16_),
	.CK(int_clk),
	.D(n1461), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__16_),
	.CK(int_clk),
	.D(n1460), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__16_),
	.CK(int_clk),
	.D(n1459), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__16_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__16_),
	.CK(int_clk),
	.D(n1458), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__17_),
	.CK(int_clk),
	.D(n1457), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__17_),
	.CK(int_clk),
	.D(n1456), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__17_),
	.CK(int_clk),
	.D(n1455), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__17_),
	.CK(int_clk),
	.D(n1454), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__17_),
	.CK(int_clk),
	.D(n1453), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__17_),
	.CK(int_clk),
	.D(n1452), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__17_),
	.CK(int_clk),
	.D(n1451), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__17_),
	.CK(int_clk),
	.D(n1449), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__17_),
	.CK(int_clk),
	.D(n1448), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__17_),
	.CK(int_clk),
	.D(n1447), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__17_),
	.CK(int_clk),
	.D(n1446), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__17_),
	.CK(int_clk),
	.D(n1445), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__17_),
	.CK(int_clk),
	.D(n1444), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__17_),
	.CK(int_clk),
	.D(n1443), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__17_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__17_),
	.CK(int_clk),
	.D(n1442), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__18_),
	.CK(int_clk),
	.D(n1441), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__18_),
	.CK(int_clk),
	.D(n1440), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__18_),
	.CK(int_clk),
	.D(n1439), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__18_),
	.CK(int_clk),
	.D(n1438), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__18_),
	.CK(int_clk),
	.D(n1437), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__18_),
	.CK(int_clk),
	.D(n1436), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__18_),
	.CK(int_clk),
	.D(n1434), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__18_),
	.CK(int_clk),
	.D(n1433), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__18_),
	.CK(int_clk),
	.D(n1432), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__18_),
	.CK(int_clk),
	.D(n1431), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__18_),
	.CK(int_clk),
	.D(n1430), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__18_),
	.CK(int_clk),
	.D(n1429), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__18_),
	.CK(int_clk),
	.D(n1428), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__18_),
	.CK(int_clk),
	.D(n1427), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__18_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__18_),
	.CK(int_clk),
	.D(n1426), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__19_),
	.CK(int_clk),
	.D(n1425), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__19_),
	.CK(int_clk),
	.D(n1424), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__19_),
	.CK(int_clk),
	.D(n1423), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__19_),
	.CK(int_clk),
	.D(n1422), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_4__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_4__19_),
	.CK(int_clk),
	.D(n1421), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__19_),
	.CK(int_clk),
	.D(n1419), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__19_),
	.CK(int_clk),
	.D(n1418), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__19_),
	.CK(int_clk),
	.D(n1417), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__19_),
	.CK(int_clk),
	.D(n1416), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__19_),
	.CK(int_clk),
	.D(n1415), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__19_),
	.CK(int_clk),
	.D(n1414), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__19_),
	.CK(int_clk),
	.D(n1413), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__19_),
	.CK(int_clk),
	.D(n1412), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__19_),
	.CK(int_clk),
	.D(n1411), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_15__19_ (
	.Q(Mfifo_psum_M_ffmem_mem_15__19_),
	.CK(int_clk),
	.D(n1410), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_0__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_0__20_),
	.CK(int_clk),
	.D(n1409), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_1__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_1__20_),
	.CK(int_clk),
	.D(n1408), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_2__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_2__20_),
	.CK(int_clk),
	.D(n1407), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_3__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_3__20_),
	.CK(int_clk),
	.D(n1406), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_5__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_5__20_),
	.CK(int_clk),
	.D(n1404), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_6__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_6__20_),
	.CK(int_clk),
	.D(n1403), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_7__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_7__20_),
	.CK(int_clk),
	.D(n1402), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_8__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_8__20_),
	.CK(int_clk),
	.D(n1401), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_9__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_9__20_),
	.CK(int_clk),
	.D(n1400), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_10__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_10__20_),
	.CK(int_clk),
	.D(n1399), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_11__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_11__20_),
	.CK(int_clk),
	.D(n1398), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_12__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_12__20_),
	.CK(int_clk),
	.D(n1397), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_13__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_13__20_),
	.CK(int_clk),
	.D(n1396), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFQX05AR9 Mfifo_psum_M_ffmem_mem_reg_14__20_ (
	.Q(Mfifo_psum_M_ffmem_mem_14__20_),
	.CK(int_clk),
	.D(n1395), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 DP_OP_1207J5_130_8771_U3 (
	.CO(DP_OP_1207J5_130_8771_n2),
	.S(C175_DATA2_4),
	.CI(DP_OP_1207J5_130_8771_n3),
	.I1(psum_addr[4]),
	.I2(Mcntl_Mcntldata_N453), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 DP_OP_1207J5_130_8771_U4 (
	.CO(DP_OP_1207J5_130_8771_n3),
	.S(C175_DATA2_3),
	.CI(DP_OP_1207J5_130_8771_n4),
	.I1(n3835),
	.I2(Mcntl_Mcntldata_N453), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX1AR9 R_21304 (
	.Q(n3830),
	.CK(int_clk),
	.D(n2076),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFSBQX1AR9 R_20585 (
	.Q(n3208),
	.CK(int_clk),
	.D(n2404),
	.SB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX8K1AR9 R_20840 (
	.Q(psum_addr[0]),
	.CK(int_clk),
	.D(n2077),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFSBQX1AR9 R_21130 (
	.Q(n3119),
	.CK(int_clk),
	.D(n2403),
	.SB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX4K1AR9 R_21190 (
	.Q(n3831),
	.CK(int_clk),
	.D(n2076),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX8K1AR9 R_21269 (
	.Q(n3841),
	.CK(int_clk),
	.D(n2076),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX8K1AR9 R_21307 (
	.Q(n3834),
	.CK(int_clk),
	.D(n2075),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX4K1AR9 R_21358 (
	.Q(psum_addr[1]),
	.CK(int_clk),
	.D(n2078),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFSBQX4K1AR9 R_21359 (
	.Q(n2912),
	.CK(int_clk),
	.D(n2401),
	.SB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX05AR9 Mcntl_Mcntldata_Mcoen_qout_r_reg_0_ (
	.Q(coen),
	.CK(int_clk),
	.D(xen4),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFSBQX1AR9 R_21306 (
	.Q(n3209),
	.CK(int_clk),
	.D(n2402),
	.SB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   DFFRBQX2AR9 Mcntl_Mcntldata_c_p_cout_reg_0_ (
	.Q(sel_ccp),
	.CK(int_clk),
	.D(n2374),
	.RB(int_rst_n), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   CLKINVX2AR9 U2524 (
	.O(n3835),
	.I(n3209), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX1AR9 U2525 (
	.O(n3842),
	.I(n3030), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X1AR9 U2526 (
	.O(adden_sec),
	.A1(n3533),
	.B1(Mcntl_Mcntldata_c_p_cin[1]),
	.B2(Mcntl_Mcntldata_c_p_cin[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2527 (
	.O(n3164),
	.I(n3090), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U2528 (
	.O(n3255),
	.A1(n3529),
	.B1(Mcntl_flag),
	.B2(n3173), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X2OAR9 U2529 (
	.O(n3821),
	.I1(n3551),
	.I2(n3553), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX1AR9 U2530 (
	.O(n2398),
	.I(n3794), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   CLKINVX2AR9 U2531 (
	.O(n3801),
	.I(n2902), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X2OAR9 U2532 (
	.O(n3799),
	.I1(n3554),
	.I2(n3553), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X2OAR9 U2533 (
	.O(n3797),
	.I1(n3552),
	.I2(n3553), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X2OAR9 U2534 (
	.O(n3813),
	.I1(n3551),
	.I2(n3545), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X2OAR9 U2535 (
	.O(n3817),
	.I1(n3545),
	.I2(n3554), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2536 (
	.O(n3252),
	.I1(n2417),
	.I2(n3080), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2537 (
	.O(n3173),
	.I1(n3080),
	.I2(n3274), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U2538 (
	.O(n3235),
	.I1(Mcntl_Mcntldata_c_x_cin[1]),
	.I2(Mcntl_Mcntldata_c_x_cin[0]),
	.I3(n3108), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND3B1X2AR9 U2539 (
	.O(n2413),
	.B3(count_k[0]),
	.I1(n3839),
	.I2(Mcntl_Mcntldata_comp_psum), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U2540 (
	.O(n2460),
	.I(n2840), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX4AR9 U2541 (
	.O(n3839),
	.I(n2412), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U2542 (
	.O(n2475),
	.I(n2869), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   CLKNAND2X1AR9 U2543 (
	.O(n3108),
	.I1(n2888),
	.I2(n3091), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX1AR9 U2544 (
	.O(n2399),
	.I(n3818), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX1AR9 U2545 (
	.O(n2400),
	.I(n3820), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2546 (
	.O(n3080),
	.I(n3532), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U2547 (
	.O(n2433),
	.I(n2860), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2548 (
	.O(n3032),
	.I1(n3030),
	.I2(n3029), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2549 (
	.O(n3529),
	.I1(Mcntl_Mcntl_current_state[0]),
	.I2(n3250), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1OAR9 U2550 (
	.O(n2861),
	.I1(Mfifo_psum_raddr[0]),
	.I2(n2440), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U2551 (
	.O(n2536),
	.I(n2825), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1OAR9 U2552 (
	.O(n2867),
	.I1(n3029),
	.I2(n2441), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U2553 (
	.O(n2614),
	.I(n2613), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U2554 (
	.O(n3558),
	.I(n3751), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2555 (
	.O(n3532),
	.I1(n3100),
	.I2(n3250), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2556 (
	.O(n3165),
	.I1(n3172),
	.I2(n3178), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X1AR9 U2557 (
	.O(n3008),
	.I1(Mfifo_coe_waddr[3]),
	.I2(n3070),
	.I3(n3012), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2558 (
	.O(n3144),
	.I1(n3224),
	.I2(n3246), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND3B2X1AR9 U2559 (
	.O(n3222),
	.B2(n3012),
	.B3(n3845),
	.I1(wen_coe_fifo), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX1AR9 U2560 (
	.O(n3030),
	.I(n2426), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U2561 (
	.O(c_k_cin[0]),
	.A1(coen),
	.A2(n2431),
	.B1B(coen),
	.B2B(Mcntl_Mcntldata_c_cin[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U2562 (
	.O(c_k_cin[1]),
	.A1(coen),
	.A2(n3111),
	.B1B(Mcntl_Mcntldata_c_cin[1]),
	.B2B(coen), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   CLKINVX8AR9 U2563 (
	.O(n3838),
	.I(n2408), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X1AR9 U2564 (
	.O(n2969),
	.I1(Mfifo_xin_waddr[3]),
	.I2(n3054),
	.I3(n2973), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U2565 (
	.O(coe_wfull),
	.I(n3845), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX1AR9 U2566 (
	.O(n3530),
	.I(Mcntl_Mcntldata_count[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX6AR9 U2567 (
	.O(n3843),
	.I(n3208), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U2568 (
	.O(psum_rempty),
	.I(n3847), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X1AR9 U2569 (
	.O(n3070),
	.B2(n3845),
	.I1(wen_coe_fifo), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X1AR9 U2570 (
	.O(n3054),
	.B2(n3846),
	.I1(wen_xin_fifo), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U2571 (
	.O(xin_wfull),
	.I(n3846), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X1AR9 U2572 (
	.O(n2426),
	.B2(n3847),
	.I1(ren_psum_fifo), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   CLKINVX2AR9 U2573 (
	.O(n3837),
	.I(n2912), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2574 (
	.O(n2401),
	.I(n2078), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX4AR9 U2575 (
	.O(n3836),
	.I(n2912), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2576 (
	.O(n2402),
	.I(n2075), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2577 (
	.O(n2404),
	.I(n2073), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2578 (
	.O(n2960),
	.I1(n2959),
	.I2(n2961), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2579 (
	.O(n2962),
	.I1(n2953),
	.I2(n2423), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2580 (
	.O(n2958),
	.I1(n2953),
	.I2(n2952), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2581 (
	.O(n2417),
	.I1(n3144),
	.I2(n3165), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 U2582 (
	.CO(DP_OP_1207J5_130_8771_n6),
	.S(C175_DATA2_0),
	.CI(DP_OP_1207J5_130_8771_n12),
	.I1(Mcntl_Mcntldata_N453),
	.I2(n3838), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2583 (
	.O(n2430),
	.I1(n3091),
	.I2(Mcntl_Mcntldata_c_W_r4[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U2584 (
	.O(n3555),
	.I1(n3549),
	.I2(Mfifo_psum_waddr[3]),
	.I3(n3548), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U2585 (
	.O(n3546),
	.I1(n3549),
	.I2(n3548),
	.I3(n3543), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2586 (
	.O(n3811),
	.I(n3780), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X1AR9 U2587 (
	.O(n2976),
	.I1(n3054),
	.I2(n3052),
	.I3(n2973), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X1AR9 U2588 (
	.O(n3015),
	.I1(n3070),
	.I2(n3068),
	.I3(n3012), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2589 (
	.O(n2888),
	.I1(Mcntl_Mcntldata_c_x_H[3]),
	.I2(n3118), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2590 (
	.O(n2425),
	.I(Mcntl_Mcntl_current_state[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X1AR9 U2591 (
	.O(n2995),
	.I1(n3052),
	.I2(n3213), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X1AR9 U2592 (
	.O(n2981),
	.I1(n3068),
	.I2(n3222), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2593 (
	.O(n2420),
	.A1(Mcntl_Mcntldata_count[1]),
	.A2(n3255),
	.B1(xen4),
	.B2(n2419), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U2594 (
	.O(n2419),
	.A1(n2418),
	.B1(c_ky[0]),
	.B2(n3087),
	.C1(n3178),
	.C2(Mcntl_Mcntldata_ky_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U2595 (
	.O(n2418),
	.A1(n3144),
	.B1(c_ky[1]),
	.B2(n3082),
	.C1(n3172),
	.C2(Mcntl_Mcntldata_ky_reg[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2596 (
	.O(n3549),
	.I1(psum_wfull),
	.I2(n3238), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2597 (
	.O(n3810),
	.I1(n3809),
	.I2(n3808),
	.I3(n3807),
	.I4(n3806), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U2598 (
	.O(n3783),
	.A1(n3782),
	.B1(n3781),
	.C1(psum2_reg3[17]),
	.C2(n2407), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U2599 (
	.O(n3733),
	.A1(n3732),
	.B1(n3731),
	.C1(psum2_reg3[9]),
	.C2(n2407), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U2600 (
	.O(n3727),
	.A1(n3726),
	.B1(n3725),
	.C1(psum1_reg3[8]),
	.C2(n3558), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U2601 (
	.O(n3715),
	.A1(n3714),
	.B1(n3713),
	.C1(n3558),
	.C2(psum1_reg3[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U2602 (
	.O(n3686),
	.A1(n3685),
	.B1(n3811),
	.B2(psum2_reg1[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U2603 (
	.O(n3680),
	.A1(n3679),
	.B1(n3678),
	.C1(n3811),
	.C2(psum2_reg1[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U2604 (
	.O(n3658),
	.A1(n3657),
	.B1(n3656),
	.C1(psum2_reg4[17]),
	.C2(n2407), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U2605 (
	.O(n3646),
	.A1(n3645),
	.B1(n3644),
	.C1(psum1_reg4[15]),
	.C2(n3558), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U2606 (
	.O(n3639),
	.A1(n3638),
	.B1(n3637),
	.C1(n3802),
	.C2(psum1_reg2[14]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U2607 (
	.O(n3581),
	.A1(n3580),
	.B1(n3579),
	.C1(psum1_reg4[4]),
	.C2(n3558), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U2608 (
	.O(n3564),
	.A1(n3563),
	.B1(n3811),
	.B2(psum2_reg2[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2609 (
	.O(n2974),
	.I1(n2993),
	.I2(n2976), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2610 (
	.O(n2977),
	.I1(n2992),
	.I2(n2976), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2611 (
	.O(n2975),
	.I1(n2994),
	.I2(n2976), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2612 (
	.O(n2978),
	.I1(n3048),
	.I2(n2976), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2613 (
	.O(n3006),
	.I1(n2995),
	.I2(n2993), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2614 (
	.O(n2996),
	.I1(n2995),
	.I2(n2992), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2615 (
	.O(n3000),
	.I1(n2995),
	.I2(n2994), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2616 (
	.O(n2967),
	.I1(n3048),
	.I2(n2969), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2617 (
	.O(n2990),
	.I1(n2989),
	.I2(n2992), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2618 (
	.O(n2991),
	.I1(n2989),
	.I2(n2994), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2619 (
	.O(n3022),
	.I1(n3013),
	.I2(n3015), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2620 (
	.O(n3018),
	.I1(n3016),
	.I2(n3015), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2621 (
	.O(n3028),
	.I1(n3014),
	.I2(n3015), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2622 (
	.O(n3024),
	.I1(n3066),
	.I2(n3015), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2623 (
	.O(n3007),
	.I1(n3066),
	.I2(n3008), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   XOR2X05AR9 U2624 (
	.O(DP_OP_1205J5_125_5849_n15),
	.I1(n2966),
	.I2(C2_Z_0), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2625 (
	.O(n2403),
	.I1(n2084),
	.I2(n2085), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2626 (
	.O(n3090),
	.I1(n3235),
	.I2(n3252), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2627 (
	.O(n3091),
	.I1(Mcntl_Mcntldata_c_W_d4[0]),
	.I2(Mcntl_Mcntldata_c_W_d4[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U2628 (
	.O(n3522),
	.I1(n3235),
	.I2(n3233),
	.I3(n3520), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 U2629 (
	.CO(n2895),
	.S(n3295),
	.CI(Mcntl_Mcntldata_ky_reg[1]),
	.I1(n3112),
	.I2(n2894), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   FAX05AR9 U2630 (
	.CO(n3187),
	.S(n3283),
	.CI(n3514),
	.I1(Mcntl_Mcntldata_kx_reg[1]),
	.I2(n3286), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2631 (
	.O(n3533),
	.I(Mcntl_Mcntldata_comp_psum), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X1AR9 U2632 (
	.O(n2412),
	.I1(n3250),
	.I2(Mcntl_Mcntldata_count[0]),
	.I3(n3530), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2633 (
	.O(n3250),
	.I1(n2425),
	.I2(Mcntl_Mcntl_current_state[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2634 (
	.O(n3246),
	.I(c_kx[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2635 (
	.O(n3224),
	.I(c_kx[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2636 (
	.O(n3274),
	.I(n2417), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2637 (
	.O(n3100),
	.I(Mcntl_Mcntl_current_state[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U2638 (
	.O(n3238),
	.I1(Mcntl_Mcntl_current_state[1]),
	.I2(Mcntl_Mcntl_current_state[2]),
	.I3(Mcntl_Mcntl_current_state[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2639 (
	.O(n3178),
	.I(c_ky[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2640 (
	.O(n3172),
	.I(c_ky[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2641 (
	.O(n3050),
	.I1(n2995),
	.I2(n3048), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX1AR9 U2642 (
	.O(n3213),
	.I(n3049), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2643 (
	.O(n3051),
	.I1(n3048),
	.I2(n2989), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2644 (
	.O(n3052),
	.I(Mfifo_xin_waddr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2645 (
	.O(n3547),
	.I1(n3193),
	.I2(n3556), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2646 (
	.O(n3037),
	.I1(n3032),
	.I2(Mfifo_psum_raddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2647 (
	.O(n3067),
	.I1(n3066),
	.I2(n2981), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2648 (
	.O(n3068),
	.I(Mfifo_coe_waddr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U2649 (
	.O(xen1),
	.B2(n3144),
	.I1(xen4), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   XNOR2X05AR9 U2650 (
	.O(n2911),
	.I1(n2910),
	.I2(psum_addr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X1AR9 U2651 (
	.O(xen4),
	.I1(n3164),
	.I2(n3173), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2652 (
	.O(n2913),
	.I(n3841), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2653 (
	.O(n2909),
	.I(n3838), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2654 (
	.O(n2920),
	.I(psum_addr[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   XOR2X05AR9 U2655 (
	.O(n3207),
	.I1(DP_OP_1205J5_125_5849_n2),
	.I2(n3204), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR4X3AR9 U2656 (
	.O(n2405),
	.I1(Mfifo_psum_raddr[0]),
	.I2(Mfifo_psum_raddr[1]),
	.I3(Mfifo_psum_raddr[3]),
	.I4(Mfifo_psum_raddr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR4X3AR9 U2657 (
	.O(n2406),
	.I1(Mfifo_psum_raddr[3]),
	.I2(Mfifo_psum_raddr[1]),
	.I3(n3029),
	.I4(n3036), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X1AR9 U2658 (
	.O(adden),
	.A1(n2420),
	.B1(Mcntl_flag),
	.B2(n3252), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X2AR9 U2659 (
	.O(n2407),
	.I1(sel_ccp),
	.I2(sel_reg[0]),
	.I3(n3537), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2660 (
	.O(Mcntl_Mcntldata_N453),
	.I1(n3147),
	.I2(n2416), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   XOR2X05AR9 U2661 (
	.O(DP_OP_1205J5_125_5849_n14),
	.I1(n2957),
	.I2(C2_Z_0), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U2662 (
	.O(n3826),
	.A1(n3810),
	.B1(n3811),
	.B2(psum2_reg1[20]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U2663 (
	.O(n3621),
	.A1(n3620),
	.B1(n3619),
	.C1(psum1_reg4[11]),
	.C2(n3751), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2664 (
	.O(n3820),
	.I1(n3551),
	.I2(n3555), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2665 (
	.O(n2988),
	.I1(n2989),
	.I2(n2993), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2666 (
	.O(n2982),
	.I1(n2981),
	.I2(n3013), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2667 (
	.O(n3027),
	.I(ext_coe[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR3B2X05AR9 U2668 (
	.O(n3267),
	.B2(n3231),
	.B3(n3104),
	.I1(coe_rempty), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2669 (
	.O(n3064),
	.I1(n3066),
	.I2(n2985), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U2670 (
	.O(n2078),
	.A1(n2925),
	.A2(n2912),
	.B1B(n2911),
	.B2B(n2923), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2671 (
	.O(Mfifo_psum_M_ffmem_N109),
	.I1(n2804),
	.I2(n2803), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2672 (
	.O(Mfifo_psum_M_ffmem_N82),
	.I1(n2674),
	.I2(n2673), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2673 (
	.O(Mfifo_psum_M_ffmem_N96),
	.I1(n2794),
	.I2(n2793), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U2674 (
	.O(n2072),
	.A1(n2919),
	.A2(n3205),
	.B1B(C174_DATA2_1),
	.B2B(n2916), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U2675 (
	.O(Mfifo_psum_M_rptr_rbinnext[2]),
	.B2(n3033),
	.I1(n3035), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX6AR9 U2676 (
	.O(n2408),
	.I(psum_addr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2677 (
	.O(n3055),
	.I(Mfifo_xin_waddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X1AR9 U2678 (
	.O(n3049),
	.I1(Mfifo_xin_waddr[0]),
	.I2(n3054), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2679 (
	.O(n3053),
	.I1(n3049),
	.I2(n3055), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA12X05AR9 U2680 (
	.O(Mfifo_xin_M_wptr_wbinnext[1]),
	.A1(n3053),
	.B1(n3055),
	.B2(n3049), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2681 (
	.O(n3544),
	.I(Mfifo_psum_waddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2682 (
	.O(n3193),
	.I1(n3549),
	.I2(Mfifo_psum_waddr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2683 (
	.O(n3194),
	.I1(n3193),
	.I2(n3544), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA12X05AR9 U2684 (
	.O(Mfifo_psum_M_wptr_wbinnext[1]),
	.A1(n3194),
	.B1(n3544),
	.B2(n3193), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2685 (
	.O(n3111),
	.I(Mcntl_Mcntldata_c_x_cin[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2686 (
	.O(n2414),
	.I1(Mcntl_Mcntldata_c_p_cout[2]),
	.I2(Mcntl_Mcntldata_c_p_cout[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2687 (
	.O(n3298),
	.I(Mcntl_Mcntldata_c_p_H[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2688 (
	.O(n3292),
	.I1(Mcntl_Mcntldata_c_p_H[0]),
	.I2(Mcntl_Mcntldata_c_p_H[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2689 (
	.O(n3303),
	.I1(n3298),
	.I2(n3292), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2690 (
	.O(n3181),
	.I1(Mcntl_Mcntldata_c_p_H[3]),
	.I2(n3303), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2691 (
	.O(n3776),
	.I1(sel_reg[1]),
	.I2(sel_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U2692 (
	.O(n3190),
	.I1(Mcntl_Mcntldata_c_p_W[2]),
	.I2(Mcntl_Mcntldata_c_p_W[3]),
	.I3(n3776), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2693 (
	.O(n3099),
	.I1(n2414),
	.I2(n3181),
	.I3(n3190),
	.I4(n3622), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2694 (
	.O(n3188),
	.I1(n3549),
	.I2(n3099), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2695 (
	.O(n3277),
	.I1(sel_ccp),
	.I2(n3188), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2696 (
	.O(n3147),
	.I1(n3277),
	.I2(n2414), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2697 (
	.O(n3640),
	.I(n3776), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2B1X05AR9 U2698 (
	.O(n2415),
	.B2(n2414),
	.I1(n3640), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U2699 (
	.O(n2907),
	.A1(n2413),
	.B1(n3277),
	.B2(n2415), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2700 (
	.O(n2416),
	.I(n2907), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2701 (
	.O(n3128),
	.I(Mcntl_Mcntldata_c_x_H[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2702 (
	.O(n3118),
	.I1(n3119),
	.I2(n3128), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2703 (
	.O(n3087),
	.I(Mcntl_Mcntldata_ky_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2704 (
	.O(n3082),
	.I(Mcntl_Mcntldata_ky_reg[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2705 (
	.O(n2915),
	.I1(xen4),
	.I2(n3246), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2706 (
	.O(n2886),
	.I1(Mcntl_Mcntldata_c_W_r4[1]),
	.I2(Mcntl_Mcntldata_c_W_r4[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2707 (
	.O(n3233),
	.I(n2886), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2708 (
	.O(n3101),
	.I(Mcntl_Mcntl_current_state[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U2709 (
	.O(n3104),
	.I1(Mcntl_Mcntl_current_state[2]),
	.I2(Mcntl_Mcntl_current_state[0]),
	.I3(n3101), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2710 (
	.O(n3232),
	.I(n3104), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2711 (
	.O(n3520),
	.I1(xin_rempty),
	.I2(n3232), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2712 (
	.O(n2914),
	.I(n3522), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI13X05AR9 U2713 (
	.O(n2421),
	.A1(n2914),
	.B1(n2915),
	.B2(n3165),
	.B3(n3108), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2714 (
	.O(n2963),
	.I1(xen1),
	.I2(n2421), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2715 (
	.O(n2422),
	.I(n2915), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2716 (
	.O(n2953),
	.I1(n2963),
	.I2(n2422), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR3X1AR9 U2717 (
	.O(n2959),
	.I1(n2953),
	.I2(n3091),
	.I3(n3165), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2B1X05AR9 U2718 (
	.O(n2423),
	.B2(n3091),
	.I1(n3165), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2719 (
	.O(n2947),
	.I(n2962), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X1AR9 U2720 (
	.O(C2_Z_0),
	.I1(n2959),
	.I2(n2947), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U2721 (
	.O(n2427),
	.I1(Mcntl_Mcntl_current_state[1]),
	.I2(Mcntl_Mcntl_current_state[2]),
	.I3(Mcntl_Mcntl_current_state[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U2722 (
	.O(int_end_send),
	.B2(int_enable),
	.I1(n2427), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2723 (
	.O(n2424),
	.I(Mcntl_Mcntldata_c_W_r4[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2724 (
	.O(n2429),
	.I(n2430), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2725 (
	.O(wen_x_reg[2]),
	.I1(n2424),
	.I2(n2429), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2726 (
	.O(wen_x_reg[0]),
	.I1(n2430),
	.I2(n2424), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U2727 (
	.O(n3228),
	.I1(count_k[0]),
	.I2(count_k[2]),
	.I3(count_k[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U2728 (
	.O(n2388),
	.A1(n3839),
	.B1(count_k[0]),
	.B2(n3228), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2729 (
	.O(n2885),
	.I1(n3100),
	.I2(Mcntl_Mcntl_current_state[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2730 (
	.O(n2883),
	.I(n2885), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2731 (
	.O(n3240),
	.I1(Mcntl_Mcntl_current_state[1]),
	.I2(n2883), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2732 (
	.O(n2428),
	.I1(n3240),
	.I2(n3104), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2733 (
	.O(Mfifo_xin_M_rptr_N1),
	.I1(xin_rempty),
	.I2(n2428), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U2734 (
	.O(n2905),
	.I1(Mcntl_Mcntl_current_state[0]),
	.I2(n2425),
	.I3(n3101), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U2735 (
	.O(int_end_comp),
	.B2(int_send),
	.I1(n2905), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U2736 (
	.O(n3829),
	.I1(n2427),
	.I2(int_enable), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   MUX2X05AR9 U2737 (
	.O(n1387),
	.I0(int_W[3]),
	.I1(Mcntl_Mcntldata_x_W_reg[3]),
	.S(n3829), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   MUX2X05AR9 U2738 (
	.O(n1388),
	.I0(int_W[2]),
	.I1(Mcntl_Mcntldata_x_W_reg[2]),
	.S(n3829), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2739 (
	.O(Mfifo_coe_M_rptr_N1),
	.I1(coe_rempty),
	.I2(n2428), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2740 (
	.O(wen_x_reg[3]),
	.I1(Mcntl_Mcntldata_c_W_r4[0]),
	.I2(n2429), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U2741 (
	.O(wen_x_reg[1]),
	.I1(Mcntl_Mcntldata_c_W_r4[0]),
	.I2(n2430), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2742 (
	.O(n2431),
	.I(Mcntl_Mcntldata_c_x_cin[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2743 (
	.O(n3029),
	.I(Mfifo_psum_raddr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U2744 (
	.O(n3031),
	.I1(Mfifo_psum_raddr[1]),
	.I2(Mfifo_psum_raddr[3]),
	.I3(Mfifo_psum_raddr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2745 (
	.O(n2825),
	.I1(n3029),
	.I2(n3031), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2746 (
	.O(n2432),
	.I(Mfifo_psum_raddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2747 (
	.O(n3036),
	.I(Mfifo_psum_raddr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U2748 (
	.O(n2442),
	.I1(Mfifo_psum_raddr[3]),
	.I2(n2432),
	.I3(n3036), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1OAR9 U2749 (
	.O(n2868),
	.I1(n3029),
	.I2(n2442), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2750 (
	.O(n2437),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__5_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR4X1AR9 U2751 (
	.O(n2872),
	.I1(Mfifo_psum_raddr[0]),
	.I2(Mfifo_psum_raddr[1]),
	.I3(Mfifo_psum_raddr[3]),
	.I4(n3036), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2752 (
	.O(n2436),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__5_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U2753 (
	.O(n2443),
	.I1(Mfifo_psum_raddr[3]),
	.I2(Mfifo_psum_raddr[2]),
	.I3(n2432), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2754 (
	.O(n2869),
	.I1(Mfifo_psum_raddr[0]),
	.I2(n2443), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2755 (
	.O(n2860),
	.I1(Mfifo_psum_raddr[0]),
	.I2(n3031), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2756 (
	.O(n2435),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__5_),
	.B1(n2433),
	.B2(Mfifo_psum_M_ffmem_mem_14__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U2757 (
	.O(n2438),
	.I1(Mfifo_psum_raddr[3]),
	.I2(Mfifo_psum_raddr[1]),
	.I3(n3036), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1OAR9 U2758 (
	.O(n2871),
	.I1(n3029),
	.I2(n2438), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2759 (
	.O(n2434),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__5_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2760 (
	.O(n2449),
	.I1(n2437),
	.I2(n2436),
	.I3(n2435),
	.I4(n2434), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U2761 (
	.O(n2439),
	.I(Mfifo_psum_raddr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U2762 (
	.O(n2441),
	.I1(Mfifo_psum_raddr[1]),
	.I2(n2439),
	.I3(n3036), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1OAR9 U2763 (
	.O(n2870),
	.I1(Mfifo_psum_raddr[0]),
	.I2(n2438), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2764 (
	.O(n2447),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__5_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U2765 (
	.O(n2440),
	.I1(Mfifo_psum_raddr[1]),
	.I2(Mfifo_psum_raddr[2]),
	.I3(n2439), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR4X1AR9 U2766 (
	.O(n2613),
	.I1(Mfifo_psum_raddr[3]),
	.I2(Mfifo_psum_raddr[1]),
	.I3(Mfifo_psum_raddr[2]),
	.I4(n3029), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2767 (
	.O(n2446),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__5_),
	.B1(n2613),
	.B2(Mfifo_psum_M_ffmem_mem_1__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U2768 (
	.O(n2840),
	.I1(n3029),
	.I2(n2440), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1OAR9 U2769 (
	.O(n2858),
	.I1(Mfifo_psum_raddr[0]),
	.I2(n2441), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2770 (
	.O(n2445),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__5_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1OAR9 U2771 (
	.O(n2862),
	.I1(Mfifo_psum_raddr[0]),
	.I2(n2442), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1OAR9 U2772 (
	.O(n2859),
	.I1(n3029),
	.I2(n2443), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2773 (
	.O(n2444),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__5_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2774 (
	.O(n2448),
	.I1(n2447),
	.I2(n2446),
	.I3(n2445),
	.I4(n2444), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2775 (
	.O(Mfifo_psum_M_ffmem_N112),
	.I1(n2449),
	.I2(n2448), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2776 (
	.O(n2453),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__34_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2777 (
	.O(n2452),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__34_),
	.B1(n2869),
	.B2(Mfifo_psum_M_ffmem_mem_12__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2778 (
	.O(n2451),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__34_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2779 (
	.O(n2450),
	.A1(n2859),
	.A2(Mfifo_psum_M_ffmem_mem_13__34_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2780 (
	.O(n2459),
	.I1(n2453),
	.I2(n2452),
	.I3(n2451),
	.I4(n2450), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2781 (
	.O(n2457),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__34_),
	.B1(n2613),
	.B2(Mfifo_psum_M_ffmem_mem_1__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2782 (
	.O(n2456),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__34_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2783 (
	.O(n2455),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__34_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2784 (
	.O(n2454),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__34_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2785 (
	.O(n2458),
	.I1(n2457),
	.I2(n2456),
	.I3(n2455),
	.I4(n2454), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2786 (
	.O(Mfifo_psum_M_ffmem_N83),
	.I1(n2459),
	.I2(n2458), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2787 (
	.O(n2464),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__10_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2788 (
	.O(n2463),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__10_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2789 (
	.O(n2462),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__10_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2790 (
	.O(n2461),
	.A1(n2433),
	.A2(Mfifo_psum_M_ffmem_mem_14__10_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2791 (
	.O(n2470),
	.I1(n2464),
	.I2(n2463),
	.I3(n2462),
	.I4(n2461), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2792 (
	.O(n2468),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__10_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2793 (
	.O(n2467),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__10_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2794 (
	.O(n2466),
	.A1(n2613),
	.A2(Mfifo_psum_M_ffmem_mem_1__10_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2795 (
	.O(n2465),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__10_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2796 (
	.O(n2469),
	.I1(n2468),
	.I2(n2467),
	.I3(n2466),
	.I4(n2465), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2797 (
	.O(Mfifo_psum_M_ffmem_N107),
	.I1(n2470),
	.I2(n2469), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2798 (
	.O(n2474),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__40_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2799 (
	.O(n2473),
	.A1(n2613),
	.A2(Mfifo_psum_M_ffmem_mem_1__40_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2800 (
	.O(n2472),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__40_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2801 (
	.O(n2471),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__40_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2802 (
	.O(n2481),
	.I1(n2474),
	.I2(n2473),
	.I3(n2472),
	.I4(n2471), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U2803 (
	.O(n2841),
	.I(n2872), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2804 (
	.O(n2479),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__40_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2805 (
	.O(n2478),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__40_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2806 (
	.O(n2477),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__40_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2807 (
	.O(n2476),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__40_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2808 (
	.O(n2480),
	.I1(n2479),
	.I2(n2478),
	.I3(n2477),
	.I4(n2476), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2809 (
	.O(Mfifo_psum_M_ffmem_N77),
	.I1(n2481),
	.I2(n2480), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2810 (
	.O(n2485),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__1_),
	.B1(n2840),
	.B2(Mfifo_psum_M_ffmem_mem_7__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2811 (
	.O(n2484),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__1_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2812 (
	.O(n2483),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__1_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2813 (
	.O(n2482),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__1_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2814 (
	.O(n2491),
	.I1(n2485),
	.I2(n2484),
	.I3(n2483),
	.I4(n2482), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2815 (
	.O(n2489),
	.A1(n2613),
	.A2(Mfifo_psum_M_ffmem_mem_1__1_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2816 (
	.O(n2488),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__1_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2817 (
	.O(n2487),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__1_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2818 (
	.O(n2486),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__1_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2819 (
	.O(n2490),
	.I1(n2489),
	.I2(n2488),
	.I3(n2487),
	.I4(n2486), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2820 (
	.O(Mfifo_psum_M_ffmem_N116),
	.I1(n2491),
	.I2(n2490), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2821 (
	.O(n2495),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__27_),
	.B1(n2613),
	.B2(Mfifo_psum_M_ffmem_mem_1__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2822 (
	.O(n2494),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__27_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2823 (
	.O(n2493),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__27_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2824 (
	.O(n2492),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__27_),
	.B1(n2840),
	.B2(Mfifo_psum_M_ffmem_mem_7__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2825 (
	.O(n2501),
	.I1(n2495),
	.I2(n2494),
	.I3(n2493),
	.I4(n2492), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2826 (
	.O(n2499),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__27_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2827 (
	.O(n2498),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__27_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2828 (
	.O(n2497),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__27_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2829 (
	.O(n2496),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__27_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2830 (
	.O(n2500),
	.I1(n2499),
	.I2(n2498),
	.I3(n2497),
	.I4(n2496), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2831 (
	.O(Mfifo_psum_M_ffmem_N90),
	.I1(n2501),
	.I2(n2500), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2832 (
	.O(n2505),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__30_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2833 (
	.O(n2504),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__30_),
	.B1(n2613),
	.B2(Mfifo_psum_M_ffmem_mem_1__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2834 (
	.O(n2503),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__30_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2835 (
	.O(n2502),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__30_),
	.B1(n2867),
	.B2(Mfifo_psum_M_ffmem_mem_3__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2836 (
	.O(n2511),
	.I1(n2505),
	.I2(n2504),
	.I3(n2503),
	.I4(n2502), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2837 (
	.O(n2509),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__30_),
	.B1(n2840),
	.B2(Mfifo_psum_M_ffmem_mem_7__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2838 (
	.O(n2508),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__30_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2839 (
	.O(n2507),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__30_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2840 (
	.O(n2506),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__30_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2841 (
	.O(n2510),
	.I1(n2509),
	.I2(n2508),
	.I3(n2507),
	.I4(n2506), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2842 (
	.O(Mfifo_psum_M_ffmem_N87),
	.I1(n2511),
	.I2(n2510), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2843 (
	.O(n2515),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__39_),
	.B1(n2613),
	.B2(Mfifo_psum_M_ffmem_mem_1__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2844 (
	.O(n2514),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__39_),
	.B1(n2840),
	.B2(Mfifo_psum_M_ffmem_mem_7__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2845 (
	.O(n2513),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__39_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2846 (
	.O(n2512),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__39_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2847 (
	.O(n2521),
	.I1(n2515),
	.I2(n2514),
	.I3(n2513),
	.I4(n2512), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2848 (
	.O(n2519),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__39_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2849 (
	.O(n2518),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__39_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2850 (
	.O(n2517),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__39_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2851 (
	.O(n2516),
	.A1(n2868),
	.A2(Mfifo_psum_M_ffmem_mem_9__39_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2852 (
	.O(n2520),
	.I1(n2519),
	.I2(n2518),
	.I3(n2517),
	.I4(n2516), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2853 (
	.O(Mfifo_psum_M_ffmem_N78),
	.I1(n2521),
	.I2(n2520), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2854 (
	.O(n2525),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__37_),
	.B1(n2613),
	.B2(Mfifo_psum_M_ffmem_mem_1__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2855 (
	.O(n2524),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__37_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2856 (
	.O(n2523),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__37_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2857 (
	.O(n2522),
	.A1(n2868),
	.A2(Mfifo_psum_M_ffmem_mem_9__37_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2858 (
	.O(n2531),
	.I1(n2525),
	.I2(n2524),
	.I3(n2523),
	.I4(n2522), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2859 (
	.O(n2529),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__37_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2860 (
	.O(n2528),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__37_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2861 (
	.O(n2527),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__37_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2862 (
	.O(n2526),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__37_),
	.B1(n2867),
	.B2(Mfifo_psum_M_ffmem_mem_3__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2863 (
	.O(n2530),
	.I1(n2529),
	.I2(n2528),
	.I3(n2527),
	.I4(n2526), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2864 (
	.O(Mfifo_psum_M_ffmem_N80),
	.I1(n2531),
	.I2(n2530), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2865 (
	.O(n2535),
	.A1(Mfifo_psum_M_ffmem_mem_13__0_),
	.A2(n2859),
	.B1(Mfifo_psum_M_ffmem_mem_1__0_),
	.B2(n2613), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2866 (
	.O(n2534),
	.A1(Mfifo_psum_M_ffmem_mem_11__0_),
	.A2(n2871),
	.B1(Mfifo_psum_M_ffmem_mem_7__0_),
	.B2(n2840), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2867 (
	.O(n2533),
	.A1(Mfifo_psum_M_ffmem_mem_2__0_),
	.A2(n2858),
	.B1(Mfifo_psum_M_ffmem_mem_10__0_),
	.B2(n2870), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2868 (
	.O(n2532),
	.A1(Mfifo_psum_M_ffmem_mem_9__0_),
	.A2(n2868),
	.B1(Mfifo_psum_M_ffmem_mem_5__0_),
	.B2(n2406), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2869 (
	.O(n2542),
	.I1(n2535),
	.I2(n2534),
	.I3(n2533),
	.I4(n2532), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2870 (
	.O(n2540),
	.A1(Mfifo_psum_M_ffmem_mem_8__0_),
	.A2(n2862),
	.B1(Mfifo_psum_M_ffmem_mem_4__0_),
	.B2(n2841), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2871 (
	.O(n2539),
	.A1(Mfifo_psum_M_ffmem_mem_15__0_),
	.A2(n2536),
	.B1(Mfifo_psum_M_ffmem_mem_3__0_),
	.B2(n2867), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2872 (
	.O(n2538),
	.A1(Mfifo_psum_M_ffmem_mem_12__0_),
	.A2(n2475),
	.B1(Mfifo_psum_M_ffmem_mem_14__0_),
	.B2(n2433), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2873 (
	.O(n2537),
	.A1(Mfifo_psum_M_ffmem_mem_0__0_),
	.A2(n2405),
	.B1(Mfifo_psum_M_ffmem_mem_6__0_),
	.B2(n2861), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2874 (
	.O(n2541),
	.I1(n2540),
	.I2(n2539),
	.I3(n2538),
	.I4(n2537), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2875 (
	.O(Mfifo_psum_M_ffmem_N117),
	.I1(n2542),
	.I2(n2541), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2876 (
	.O(n2546),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__32_),
	.B1(n2840),
	.B2(Mfifo_psum_M_ffmem_mem_7__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2877 (
	.O(n2545),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__32_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2878 (
	.O(n2544),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__32_),
	.B1(n2613),
	.B2(Mfifo_psum_M_ffmem_mem_1__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2879 (
	.O(n2543),
	.A1(n2858),
	.A2(Mfifo_psum_M_ffmem_mem_2__32_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2880 (
	.O(n2552),
	.I1(n2546),
	.I2(n2545),
	.I3(n2544),
	.I4(n2543), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2881 (
	.O(n2550),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__32_),
	.B1(n2862),
	.B2(Mfifo_psum_M_ffmem_mem_8__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2882 (
	.O(n2549),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__32_),
	.B1(n2869),
	.B2(Mfifo_psum_M_ffmem_mem_12__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2883 (
	.O(n2548),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__32_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2884 (
	.O(n2547),
	.A1(n2433),
	.A2(Mfifo_psum_M_ffmem_mem_14__32_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2885 (
	.O(n2551),
	.I1(n2550),
	.I2(n2549),
	.I3(n2548),
	.I4(n2547), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2886 (
	.O(Mfifo_psum_M_ffmem_N85),
	.I1(n2552),
	.I2(n2551), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2887 (
	.O(n2556),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__3_),
	.B1(n2841),
	.B2(Mfifo_psum_M_ffmem_mem_4__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2888 (
	.O(n2555),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__3_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2889 (
	.O(n2554),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__3_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2890 (
	.O(n2553),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__3_),
	.B1(n2613),
	.B2(Mfifo_psum_M_ffmem_mem_1__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2891 (
	.O(n2562),
	.I1(n2556),
	.I2(n2555),
	.I3(n2554),
	.I4(n2553), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2892 (
	.O(n2560),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__3_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2893 (
	.O(n2559),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__3_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2894 (
	.O(n2558),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__3_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2895 (
	.O(n2557),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__3_),
	.B1(n2433),
	.B2(Mfifo_psum_M_ffmem_mem_14__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2896 (
	.O(n2561),
	.I1(n2560),
	.I2(n2559),
	.I3(n2558),
	.I4(n2557), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2897 (
	.O(Mfifo_psum_M_ffmem_N114),
	.I1(n2562),
	.I2(n2561), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2898 (
	.O(n2566),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__33_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2899 (
	.O(n2565),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__33_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2900 (
	.O(n2564),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__33_),
	.B1(n2841),
	.B2(Mfifo_psum_M_ffmem_mem_4__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2901 (
	.O(n2563),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__33_),
	.B1(n2613),
	.B2(Mfifo_psum_M_ffmem_mem_1__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2902 (
	.O(n2572),
	.I1(n2566),
	.I2(n2565),
	.I3(n2564),
	.I4(n2563), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2903 (
	.O(n2570),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__33_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2904 (
	.O(n2569),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__33_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2905 (
	.O(n2568),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__33_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2906 (
	.O(n2567),
	.A1(n2868),
	.A2(Mfifo_psum_M_ffmem_mem_9__33_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2907 (
	.O(n2571),
	.I1(n2570),
	.I2(n2569),
	.I3(n2568),
	.I4(n2567), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2908 (
	.O(Mfifo_psum_M_ffmem_N84),
	.I1(n2572),
	.I2(n2571), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2909 (
	.O(n2576),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__29_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2910 (
	.O(n2575),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__29_),
	.B1(n2841),
	.B2(Mfifo_psum_M_ffmem_mem_4__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2911 (
	.O(n2574),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__29_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2912 (
	.O(n2573),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__29_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2913 (
	.O(n2582),
	.I1(n2576),
	.I2(n2575),
	.I3(n2574),
	.I4(n2573), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2914 (
	.O(n2580),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__29_),
	.B1(n2613),
	.B2(Mfifo_psum_M_ffmem_mem_1__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2915 (
	.O(n2579),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__29_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2916 (
	.O(n2578),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__29_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2917 (
	.O(n2577),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__29_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2918 (
	.O(n2581),
	.I1(n2580),
	.I2(n2579),
	.I3(n2578),
	.I4(n2577), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2919 (
	.O(Mfifo_psum_M_ffmem_N88),
	.I1(n2582),
	.I2(n2581), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2920 (
	.O(n2586),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__22_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2921 (
	.O(n2585),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__22_),
	.B1(n2841),
	.B2(Mfifo_psum_M_ffmem_mem_4__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2922 (
	.O(n2584),
	.A1(n2433),
	.A2(Mfifo_psum_M_ffmem_mem_14__22_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2923 (
	.O(n2583),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__22_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2924 (
	.O(n2592),
	.I1(n2586),
	.I2(n2585),
	.I3(n2584),
	.I4(n2583), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2925 (
	.O(n2590),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__22_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2926 (
	.O(n2589),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__22_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2927 (
	.O(n2588),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__22_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2928 (
	.O(n2587),
	.A1(n2613),
	.A2(Mfifo_psum_M_ffmem_mem_1__22_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2929 (
	.O(n2591),
	.I1(n2590),
	.I2(n2589),
	.I3(n2588),
	.I4(n2587), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2930 (
	.O(Mfifo_psum_M_ffmem_N95),
	.I1(n2592),
	.I2(n2591), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2931 (
	.O(n2596),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__12_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2932 (
	.O(n2595),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__12_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2933 (
	.O(n2594),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__12_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2934 (
	.O(n2593),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__12_),
	.B1(n2841),
	.B2(Mfifo_psum_M_ffmem_mem_4__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2935 (
	.O(n2602),
	.I1(n2596),
	.I2(n2595),
	.I3(n2594),
	.I4(n2593), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2936 (
	.O(n2600),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__12_),
	.B1(n2433),
	.B2(Mfifo_psum_M_ffmem_mem_14__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2937 (
	.O(n2599),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__12_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2938 (
	.O(n2598),
	.A1(n2613),
	.A2(Mfifo_psum_M_ffmem_mem_1__12_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2939 (
	.O(n2597),
	.A1(n2859),
	.A2(Mfifo_psum_M_ffmem_mem_13__12_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2940 (
	.O(n2601),
	.I1(n2600),
	.I2(n2599),
	.I3(n2598),
	.I4(n2597), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2941 (
	.O(Mfifo_psum_M_ffmem_N105),
	.I1(n2602),
	.I2(n2601), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2942 (
	.O(n2606),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__2_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2943 (
	.O(n2605),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__2_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2944 (
	.O(n2604),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__2_),
	.B1(n2613),
	.B2(Mfifo_psum_M_ffmem_mem_1__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2945 (
	.O(n2603),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__2_),
	.B1(n2841),
	.B2(Mfifo_psum_M_ffmem_mem_4__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2946 (
	.O(n2612),
	.I1(n2606),
	.I2(n2605),
	.I3(n2604),
	.I4(n2603), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2947 (
	.O(n2610),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__2_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2948 (
	.O(n2609),
	.A1(n2406),
	.A2(Mfifo_psum_M_ffmem_mem_5__2_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2949 (
	.O(n2608),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__2_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2950 (
	.O(n2607),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__2_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2951 (
	.O(n2611),
	.I1(n2610),
	.I2(n2609),
	.I3(n2608),
	.I4(n2607), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2952 (
	.O(Mfifo_psum_M_ffmem_N115),
	.I1(n2612),
	.I2(n2611), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2953 (
	.O(n2618),
	.A1(n2614),
	.A2(Mfifo_psum_M_ffmem_mem_1__11_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2954 (
	.O(n2617),
	.A1(n2858),
	.A2(Mfifo_psum_M_ffmem_mem_2__11_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2955 (
	.O(n2616),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__11_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2956 (
	.O(n2615),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__11_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2957 (
	.O(n2624),
	.I1(n2618),
	.I2(n2617),
	.I3(n2616),
	.I4(n2615), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2958 (
	.O(n2622),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__11_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2959 (
	.O(n2621),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__11_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2960 (
	.O(n2620),
	.A1(n2475),
	.A2(Mfifo_psum_M_ffmem_mem_12__11_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2961 (
	.O(n2619),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__11_),
	.B1(n2433),
	.B2(Mfifo_psum_M_ffmem_mem_14__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2962 (
	.O(n2623),
	.I1(n2622),
	.I2(n2621),
	.I3(n2620),
	.I4(n2619), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2963 (
	.O(Mfifo_psum_M_ffmem_N106),
	.I1(n2624),
	.I2(n2623), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2964 (
	.O(n2628),
	.A1(n2614),
	.A2(Mfifo_psum_M_ffmem_mem_1__41_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2965 (
	.O(n2627),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__41_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2966 (
	.O(n2626),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__41_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2967 (
	.O(n2625),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__41_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2968 (
	.O(n2634),
	.I1(n2628),
	.I2(n2627),
	.I3(n2626),
	.I4(n2625), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2969 (
	.O(n2632),
	.A1(n2858),
	.A2(Mfifo_psum_M_ffmem_mem_2__41_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2970 (
	.O(n2631),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__41_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2971 (
	.O(n2630),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__41_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2972 (
	.O(n2629),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__41_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2973 (
	.O(n2633),
	.I1(n2632),
	.I2(n2631),
	.I3(n2630),
	.I4(n2629), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2974 (
	.O(Mfifo_psum_M_ffmem_N76),
	.I1(n2634),
	.I2(n2633), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2975 (
	.O(n2638),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__13_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2976 (
	.O(n2637),
	.A1(n2614),
	.A2(Mfifo_psum_M_ffmem_mem_1__13_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2977 (
	.O(n2636),
	.A1(n2433),
	.A2(Mfifo_psum_M_ffmem_mem_14__13_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2978 (
	.O(n2635),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__13_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2979 (
	.O(n2644),
	.I1(n2638),
	.I2(n2637),
	.I3(n2636),
	.I4(n2635), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2980 (
	.O(n2642),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__13_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2981 (
	.O(n2641),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__13_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2982 (
	.O(n2640),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__13_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2983 (
	.O(n2639),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__13_),
	.B1(n2862),
	.B2(Mfifo_psum_M_ffmem_mem_8__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2984 (
	.O(n2643),
	.I1(n2642),
	.I2(n2641),
	.I3(n2640),
	.I4(n2639), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2985 (
	.O(Mfifo_psum_M_ffmem_N104),
	.I1(n2644),
	.I2(n2643), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2986 (
	.O(n2648),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__7_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2987 (
	.O(n2647),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__7_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2988 (
	.O(n2646),
	.A1(n2614),
	.A2(Mfifo_psum_M_ffmem_mem_1__7_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2989 (
	.O(n2645),
	.A1(n2859),
	.A2(Mfifo_psum_M_ffmem_mem_13__7_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2990 (
	.O(n2654),
	.I1(n2648),
	.I2(n2647),
	.I3(n2646),
	.I4(n2645), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2991 (
	.O(n2652),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__7_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2992 (
	.O(n2651),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__7_),
	.B1(n2433),
	.B2(Mfifo_psum_M_ffmem_mem_14__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2993 (
	.O(n2650),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__7_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2994 (
	.O(n2649),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__7_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U2995 (
	.O(n2653),
	.I1(n2652),
	.I2(n2651),
	.I3(n2650),
	.I4(n2649), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U2996 (
	.O(Mfifo_psum_M_ffmem_N110),
	.I1(n2654),
	.I2(n2653), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2997 (
	.O(n2658),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__24_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2998 (
	.O(n2657),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__24_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U2999 (
	.O(n2656),
	.A1(n2614),
	.A2(Mfifo_psum_M_ffmem_mem_1__24_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3000 (
	.O(n2655),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__24_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3001 (
	.O(n2664),
	.I1(n2658),
	.I2(n2657),
	.I3(n2656),
	.I4(n2655), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3002 (
	.O(n2662),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__24_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3003 (
	.O(n2661),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__24_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3004 (
	.O(n2660),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__24_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3005 (
	.O(n2659),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__24_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3006 (
	.O(n2663),
	.I1(n2662),
	.I2(n2661),
	.I3(n2660),
	.I4(n2659), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3007 (
	.O(Mfifo_psum_M_ffmem_N93),
	.I1(n2664),
	.I2(n2663), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3008 (
	.O(n2668),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__35_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3009 (
	.O(n2667),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__35_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3010 (
	.O(n2666),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__35_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3011 (
	.O(n2665),
	.A1(n2614),
	.A2(Mfifo_psum_M_ffmem_mem_1__35_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3012 (
	.O(n2674),
	.I1(n2668),
	.I2(n2667),
	.I3(n2666),
	.I4(n2665), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3013 (
	.O(n2672),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__35_),
	.B1(n2840),
	.B2(Mfifo_psum_M_ffmem_mem_7__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3014 (
	.O(n2671),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__35_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3015 (
	.O(n2670),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__35_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3016 (
	.O(n2669),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__35_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3017 (
	.O(n2673),
	.I1(n2672),
	.I2(n2671),
	.I3(n2670),
	.I4(n2669), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3018 (
	.O(n2678),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__4_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3019 (
	.O(n2677),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__4_),
	.B1(n2433),
	.B2(Mfifo_psum_M_ffmem_mem_14__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3020 (
	.O(n2676),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__4_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3021 (
	.O(n2675),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__4_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3022 (
	.O(n2684),
	.I1(n2678),
	.I2(n2677),
	.I3(n2676),
	.I4(n2675), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3023 (
	.O(n2682),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__4_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3024 (
	.O(n2681),
	.A1(n2406),
	.A2(Mfifo_psum_M_ffmem_mem_5__4_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3025 (
	.O(n2680),
	.A1(n2614),
	.A2(Mfifo_psum_M_ffmem_mem_1__4_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3026 (
	.O(n2679),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__4_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3027 (
	.O(n2683),
	.I1(n2682),
	.I2(n2681),
	.I3(n2680),
	.I4(n2679), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3028 (
	.O(Mfifo_psum_M_ffmem_N113),
	.I1(n2684),
	.I2(n2683), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3029 (
	.O(n2688),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__6_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3030 (
	.O(n2687),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__6_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3031 (
	.O(n2686),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__6_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3032 (
	.O(n2685),
	.A1(n2868),
	.A2(Mfifo_psum_M_ffmem_mem_9__6_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3033 (
	.O(n2694),
	.I1(n2688),
	.I2(n2687),
	.I3(n2686),
	.I4(n2685), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3034 (
	.O(n2692),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__6_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3035 (
	.O(n2691),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__6_),
	.B1(n2862),
	.B2(Mfifo_psum_M_ffmem_mem_8__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3036 (
	.O(n2690),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__6_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3037 (
	.O(n2689),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__6_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3038 (
	.O(n2693),
	.I1(n2692),
	.I2(n2691),
	.I3(n2690),
	.I4(n2689), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3039 (
	.O(Mfifo_psum_M_ffmem_N111),
	.I1(n2694),
	.I2(n2693), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3040 (
	.O(n2698),
	.A1(n2859),
	.A2(Mfifo_psum_M_ffmem_mem_13__9_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3041 (
	.O(n2697),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__9_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3042 (
	.O(n2696),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__9_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3043 (
	.O(n2695),
	.A1(n2868),
	.A2(Mfifo_psum_M_ffmem_mem_9__9_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3044 (
	.O(n2704),
	.I1(n2698),
	.I2(n2697),
	.I3(n2696),
	.I4(n2695), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3045 (
	.O(n2702),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__9_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3046 (
	.O(n2701),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__9_),
	.B1(n2433),
	.B2(Mfifo_psum_M_ffmem_mem_14__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3047 (
	.O(n2700),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__9_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3048 (
	.O(n2699),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__9_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3049 (
	.O(n2703),
	.I1(n2702),
	.I2(n2701),
	.I3(n2700),
	.I4(n2699), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3050 (
	.O(Mfifo_psum_M_ffmem_N108),
	.I1(n2704),
	.I2(n2703), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3051 (
	.O(n2708),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__14_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3052 (
	.O(n2707),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__14_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3053 (
	.O(n2706),
	.A1(n2868),
	.A2(Mfifo_psum_M_ffmem_mem_9__14_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3054 (
	.O(n2705),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__14_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3055 (
	.O(n2714),
	.I1(n2708),
	.I2(n2707),
	.I3(n2706),
	.I4(n2705), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3056 (
	.O(n2712),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__14_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3057 (
	.O(n2711),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__14_),
	.B1(n2841),
	.B2(Mfifo_psum_M_ffmem_mem_4__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3058 (
	.O(n2710),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__14_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3059 (
	.O(n2709),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__14_),
	.B1(n2433),
	.B2(Mfifo_psum_M_ffmem_mem_14__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3060 (
	.O(n2713),
	.I1(n2712),
	.I2(n2711),
	.I3(n2710),
	.I4(n2709), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3061 (
	.O(Mfifo_psum_M_ffmem_N103),
	.I1(n2714),
	.I2(n2713), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3062 (
	.O(n2718),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__23_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3063 (
	.O(n2717),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__23_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3064 (
	.O(n2716),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__23_),
	.B1(n2840),
	.B2(Mfifo_psum_M_ffmem_mem_7__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3065 (
	.O(n2715),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__23_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3066 (
	.O(n2724),
	.I1(n2718),
	.I2(n2717),
	.I3(n2716),
	.I4(n2715), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3067 (
	.O(n2722),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__23_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3068 (
	.O(n2721),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__23_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3069 (
	.O(n2720),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__23_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3070 (
	.O(n2719),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__23_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3071 (
	.O(n2723),
	.I1(n2722),
	.I2(n2721),
	.I3(n2720),
	.I4(n2719), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3072 (
	.O(Mfifo_psum_M_ffmem_N94),
	.I1(n2724),
	.I2(n2723), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3073 (
	.O(n2728),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__36_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3074 (
	.O(n2727),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__36_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3075 (
	.O(n2726),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__36_),
	.B1(n2840),
	.B2(Mfifo_psum_M_ffmem_mem_7__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3076 (
	.O(n2725),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__36_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3077 (
	.O(n2734),
	.I1(n2728),
	.I2(n2727),
	.I3(n2726),
	.I4(n2725), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3078 (
	.O(n2732),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__36_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3079 (
	.O(n2731),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__36_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3080 (
	.O(n2730),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__36_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3081 (
	.O(n2729),
	.A1(n2858),
	.A2(Mfifo_psum_M_ffmem_mem_2__36_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3082 (
	.O(n2733),
	.I1(n2732),
	.I2(n2731),
	.I3(n2730),
	.I4(n2729), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3083 (
	.O(Mfifo_psum_M_ffmem_N81),
	.I1(n2734),
	.I2(n2733), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3084 (
	.O(n2738),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__16_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3085 (
	.O(n2737),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__16_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3086 (
	.O(n2736),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__16_),
	.B1(n2869),
	.B2(Mfifo_psum_M_ffmem_mem_12__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3087 (
	.O(n2735),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__16_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3088 (
	.O(n2744),
	.I1(n2738),
	.I2(n2737),
	.I3(n2736),
	.I4(n2735), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3089 (
	.O(n2742),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__16_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3090 (
	.O(n2741),
	.A1(n2433),
	.A2(Mfifo_psum_M_ffmem_mem_14__16_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3091 (
	.O(n2740),
	.A1(n2406),
	.A2(Mfifo_psum_M_ffmem_mem_5__16_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3092 (
	.O(n2739),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__16_),
	.B1(n2867),
	.B2(Mfifo_psum_M_ffmem_mem_3__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3093 (
	.O(n2743),
	.I1(n2742),
	.I2(n2741),
	.I3(n2740),
	.I4(n2739), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3094 (
	.O(Mfifo_psum_M_ffmem_N101),
	.I1(n2744),
	.I2(n2743), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3095 (
	.O(n2748),
	.A1(n2859),
	.A2(Mfifo_psum_M_ffmem_mem_13__31_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3096 (
	.O(n2747),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__31_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3097 (
	.O(n2746),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__31_),
	.B1(n2840),
	.B2(Mfifo_psum_M_ffmem_mem_7__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3098 (
	.O(n2745),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__31_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3099 (
	.O(n2754),
	.I1(n2748),
	.I2(n2747),
	.I3(n2746),
	.I4(n2745), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3100 (
	.O(n2752),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__31_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3101 (
	.O(n2751),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__31_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3102 (
	.O(n2750),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__31_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3103 (
	.O(n2749),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__31_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3104 (
	.O(n2753),
	.I1(n2752),
	.I2(n2751),
	.I3(n2750),
	.I4(n2749), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3105 (
	.O(Mfifo_psum_M_ffmem_N86),
	.I1(n2754),
	.I2(n2753), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3106 (
	.O(n2758),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__17_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3107 (
	.O(n2757),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__17_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3108 (
	.O(n2756),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__17_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3109 (
	.O(n2755),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__17_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3110 (
	.O(n2764),
	.I1(n2758),
	.I2(n2757),
	.I3(n2756),
	.I4(n2755), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3111 (
	.O(n2762),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__17_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3112 (
	.O(n2761),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__17_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3113 (
	.O(n2760),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__17_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3114 (
	.O(n2759),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__17_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3115 (
	.O(n2763),
	.I1(n2762),
	.I2(n2761),
	.I3(n2760),
	.I4(n2759), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3116 (
	.O(Mfifo_psum_M_ffmem_N100),
	.I1(n2764),
	.I2(n2763), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3117 (
	.O(n2768),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__20_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3118 (
	.O(n2767),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__20_),
	.B1(n2867),
	.B2(Mfifo_psum_M_ffmem_mem_3__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3119 (
	.O(n2766),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__20_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3120 (
	.O(n2765),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__20_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3121 (
	.O(n2774),
	.I1(n2768),
	.I2(n2767),
	.I3(n2766),
	.I4(n2765), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3122 (
	.O(n2772),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__20_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3123 (
	.O(n2771),
	.A1(n2460),
	.A2(Mfifo_psum_M_ffmem_mem_7__20_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3124 (
	.O(n2770),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__20_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3125 (
	.O(n2769),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__20_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3126 (
	.O(n2773),
	.I1(n2772),
	.I2(n2771),
	.I3(n2770),
	.I4(n2769), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3127 (
	.O(Mfifo_psum_M_ffmem_N97),
	.I1(n2774),
	.I2(n2773), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3128 (
	.O(n2778),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__28_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3129 (
	.O(n2777),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__28_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3130 (
	.O(n2776),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__28_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3131 (
	.O(n2775),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__28_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3132 (
	.O(n2784),
	.I1(n2778),
	.I2(n2777),
	.I3(n2776),
	.I4(n2775), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3133 (
	.O(n2782),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__28_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3134 (
	.O(n2781),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__28_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3135 (
	.O(n2780),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__28_),
	.B1(n2869),
	.B2(Mfifo_psum_M_ffmem_mem_12__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3136 (
	.O(n2779),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__28_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3137 (
	.O(n2783),
	.I1(n2782),
	.I2(n2781),
	.I3(n2780),
	.I4(n2779), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3138 (
	.O(Mfifo_psum_M_ffmem_N89),
	.I1(n2784),
	.I2(n2783), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3139 (
	.O(n2788),
	.A1(n2840),
	.A2(Mfifo_psum_M_ffmem_mem_7__21_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3140 (
	.O(n2787),
	.A1(n2859),
	.A2(Mfifo_psum_M_ffmem_mem_13__21_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3141 (
	.O(n2786),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__21_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3142 (
	.O(n2785),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__21_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3143 (
	.O(n2794),
	.I1(n2788),
	.I2(n2787),
	.I3(n2786),
	.I4(n2785), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3144 (
	.O(n2792),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__21_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3145 (
	.O(n2791),
	.A1(n2868),
	.A2(Mfifo_psum_M_ffmem_mem_9__21_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3146 (
	.O(n2790),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__21_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3147 (
	.O(n2789),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__21_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3148 (
	.O(n2793),
	.I1(n2792),
	.I2(n2791),
	.I3(n2790),
	.I4(n2789), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3149 (
	.O(n2798),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__8_),
	.B1(n2862),
	.B2(Mfifo_psum_M_ffmem_mem_8__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3150 (
	.O(n2797),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__8_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3151 (
	.O(n2796),
	.A1(n2868),
	.A2(Mfifo_psum_M_ffmem_mem_9__8_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3152 (
	.O(n2795),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__8_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3153 (
	.O(n2804),
	.I1(n2798),
	.I2(n2797),
	.I3(n2796),
	.I4(n2795), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3154 (
	.O(n2802),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__8_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3155 (
	.O(n2801),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__8_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3156 (
	.O(n2800),
	.A1(n2859),
	.A2(Mfifo_psum_M_ffmem_mem_13__8_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3157 (
	.O(n2799),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__8_),
	.B1(n2433),
	.B2(Mfifo_psum_M_ffmem_mem_14__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3158 (
	.O(n2803),
	.I1(n2802),
	.I2(n2801),
	.I3(n2800),
	.I4(n2799), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3159 (
	.O(n2808),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__15_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3160 (
	.O(n2807),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__15_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3161 (
	.O(n2806),
	.A1(n2868),
	.A2(Mfifo_psum_M_ffmem_mem_9__15_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3162 (
	.O(n2805),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__15_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3163 (
	.O(n2814),
	.I1(n2808),
	.I2(n2807),
	.I3(n2806),
	.I4(n2805), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3164 (
	.O(n2812),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__15_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3165 (
	.O(n2811),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__15_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3166 (
	.O(n2810),
	.A1(n2460),
	.A2(Mfifo_psum_M_ffmem_mem_7__15_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3167 (
	.O(n2809),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__15_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3168 (
	.O(n2813),
	.I1(n2812),
	.I2(n2811),
	.I3(n2810),
	.I4(n2809), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3169 (
	.O(Mfifo_psum_M_ffmem_N102),
	.I1(n2814),
	.I2(n2813), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3170 (
	.O(n2818),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__38_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3171 (
	.O(n2817),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__38_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3172 (
	.O(n2816),
	.A1(n2868),
	.A2(Mfifo_psum_M_ffmem_mem_9__38_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3173 (
	.O(n2815),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__38_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3174 (
	.O(n2824),
	.I1(n2818),
	.I2(n2817),
	.I3(n2816),
	.I4(n2815), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3175 (
	.O(n2822),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__38_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3176 (
	.O(n2821),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__38_),
	.B1(n2840),
	.B2(Mfifo_psum_M_ffmem_mem_7__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3177 (
	.O(n2820),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__38_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3178 (
	.O(n2819),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__38_),
	.B1(n2861),
	.B2(Mfifo_psum_M_ffmem_mem_6__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3179 (
	.O(n2823),
	.I1(n2822),
	.I2(n2821),
	.I3(n2820),
	.I4(n2819), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3180 (
	.O(Mfifo_psum_M_ffmem_N79),
	.I1(n2824),
	.I2(n2823), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3181 (
	.O(n2829),
	.A1(n2859),
	.A2(Mfifo_psum_M_ffmem_mem_13__26_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3182 (
	.O(n2828),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__26_),
	.B1(n2405),
	.B2(Mfifo_psum_M_ffmem_mem_0__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3183 (
	.O(n2827),
	.A1(n2825),
	.A2(Mfifo_psum_M_ffmem_mem_15__26_),
	.B1(n2475),
	.B2(Mfifo_psum_M_ffmem_mem_12__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3184 (
	.O(n2826),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__26_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3185 (
	.O(n2835),
	.I1(n2829),
	.I2(n2828),
	.I3(n2827),
	.I4(n2826), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3186 (
	.O(n2833),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__26_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3187 (
	.O(n2832),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__26_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3188 (
	.O(n2831),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__26_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3189 (
	.O(n2830),
	.A1(n2460),
	.A2(Mfifo_psum_M_ffmem_mem_7__26_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3190 (
	.O(n2834),
	.I1(n2833),
	.I2(n2832),
	.I3(n2831),
	.I4(n2830), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3191 (
	.O(Mfifo_psum_M_ffmem_N91),
	.I1(n2835),
	.I2(n2834), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3192 (
	.O(n2839),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__25_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3193 (
	.O(n2838),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__25_),
	.B1(n2862),
	.B2(Mfifo_psum_M_ffmem_mem_8__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3194 (
	.O(n2837),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__25_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3195 (
	.O(n2836),
	.A1(n2868),
	.A2(Mfifo_psum_M_ffmem_mem_9__25_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3196 (
	.O(n2847),
	.I1(n2839),
	.I2(n2838),
	.I3(n2837),
	.I4(n2836), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3197 (
	.O(n2845),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__25_),
	.B1(n2840),
	.B2(Mfifo_psum_M_ffmem_mem_7__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3198 (
	.O(n2844),
	.A1(n2841),
	.A2(Mfifo_psum_M_ffmem_mem_4__25_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3199 (
	.O(n2843),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__25_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3200 (
	.O(n2842),
	.A1(n2860),
	.A2(Mfifo_psum_M_ffmem_mem_14__25_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3201 (
	.O(n2846),
	.I1(n2845),
	.I2(n2844),
	.I3(n2843),
	.I4(n2842), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3202 (
	.O(Mfifo_psum_M_ffmem_N92),
	.I1(n2847),
	.I2(n2846), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3203 (
	.O(n2851),
	.A1(n2406),
	.A2(Mfifo_psum_M_ffmem_mem_5__18_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3204 (
	.O(n2850),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__18_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3205 (
	.O(n2849),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__18_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3206 (
	.O(n2848),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__18_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3207 (
	.O(n2857),
	.I1(n2851),
	.I2(n2850),
	.I3(n2849),
	.I4(n2848), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3208 (
	.O(n2855),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__18_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3209 (
	.O(n2854),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__18_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3210 (
	.O(n2853),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__18_),
	.B1(n2871),
	.B2(Mfifo_psum_M_ffmem_mem_11__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3211 (
	.O(n2852),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__18_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3212 (
	.O(n2856),
	.I1(n2855),
	.I2(n2854),
	.I3(n2853),
	.I4(n2852), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3213 (
	.O(Mfifo_psum_M_ffmem_N99),
	.I1(n2857),
	.I2(n2856), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3214 (
	.O(n2866),
	.A1(n2405),
	.A2(Mfifo_psum_M_ffmem_mem_0__19_),
	.B1(n2858),
	.B2(Mfifo_psum_M_ffmem_mem_2__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3215 (
	.O(n2865),
	.A1(n2536),
	.A2(Mfifo_psum_M_ffmem_mem_15__19_),
	.B1(n2859),
	.B2(Mfifo_psum_M_ffmem_mem_13__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3216 (
	.O(n2864),
	.A1(n2861),
	.A2(Mfifo_psum_M_ffmem_mem_6__19_),
	.B1(n2860),
	.B2(Mfifo_psum_M_ffmem_mem_14__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3217 (
	.O(n2863),
	.A1(n2862),
	.A2(Mfifo_psum_M_ffmem_mem_8__19_),
	.B1(n2460),
	.B2(Mfifo_psum_M_ffmem_mem_7__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3218 (
	.O(n2878),
	.I1(n2866),
	.I2(n2865),
	.I3(n2864),
	.I4(n2863), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3219 (
	.O(n2876),
	.A1(n2867),
	.A2(Mfifo_psum_M_ffmem_mem_3__19_),
	.B1(n2406),
	.B2(Mfifo_psum_M_ffmem_mem_5__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3220 (
	.O(n2875),
	.A1(n2869),
	.A2(Mfifo_psum_M_ffmem_mem_12__19_),
	.B1(n2868),
	.B2(Mfifo_psum_M_ffmem_mem_9__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3221 (
	.O(n2874),
	.A1(n2871),
	.A2(Mfifo_psum_M_ffmem_mem_11__19_),
	.B1(n2870),
	.B2(Mfifo_psum_M_ffmem_mem_10__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3222 (
	.O(n2873),
	.A1(n2872),
	.A2(Mfifo_psum_M_ffmem_mem_4__19_),
	.B1(n2614),
	.B2(Mfifo_psum_M_ffmem_mem_1__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3223 (
	.O(n2877),
	.I1(n2876),
	.I2(n2875),
	.I3(n2874),
	.I4(n2873), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2X05AR9 U3224 (
	.O(Mfifo_psum_M_ffmem_N98),
	.I1(n2878),
	.I2(n2877), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3225 (
	.O(n3012),
	.I(Mfifo_coe_waddr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3226 (
	.O(n3065),
	.I(n3222), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3227 (
	.O(n3071),
	.I(Mfifo_coe_waddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3228 (
	.O(n3069),
	.I1(n3071),
	.I2(n3065), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA12X05AR9 U3229 (
	.O(Mfifo_coe_M_wptr_wbinnext[1]),
	.A1(n3069),
	.B1(n3065),
	.B2(n3071), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3230 (
	.O(n2879),
	.I1(n3032),
	.I2(Mfifo_psum_raddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3231 (
	.O(n3035),
	.I1(n2879),
	.I2(n3036), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3232 (
	.O(n3033),
	.I1(n2879),
	.I2(n3036), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3233 (
	.O(n3827),
	.I(n3829), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA22X05AR9 U3234 (
	.O(n1383),
	.A1(n3827),
	.A2(Mcntl_Mcntldata_x_H_reg[3]),
	.B1(n3829),
	.B2(int_H[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA22X05AR9 U3235 (
	.O(n1384),
	.A1(n3827),
	.A2(Mcntl_Mcntldata_x_H_reg[2]),
	.B1(n3829),
	.B2(int_H[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA22X05AR9 U3236 (
	.O(n1385),
	.A1(n3827),
	.A2(Mcntl_Mcntldata_x_H_reg[1]),
	.B1(n3829),
	.B2(int_H[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3237 (
	.O(n3418),
	.I(Mfifo_xin_raddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3238 (
	.O(n2882),
	.I1(Mfifo_xin_M_rptr_N1),
	.I2(Mfifo_xin_raddr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3239 (
	.O(n3133),
	.I1(n3418),
	.I2(n2882), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3240 (
	.O(n2880),
	.I1(n3418),
	.I2(n2882), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U3241 (
	.O(Mfifo_xin_M_rptr_rbinnext[1]),
	.B2(n2880),
	.I1(n3133), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3242 (
	.O(n2881),
	.I1(Mfifo_xin_raddr[2]),
	.I2(n2880), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3243 (
	.O(n3132),
	.I1(Mfifo_xin_raddr[2]),
	.I2(n2880), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U3244 (
	.O(Mfifo_xin_M_rptr_rbinnext[2]),
	.B2(n3132),
	.I1(n2881), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3245 (
	.O(n3419),
	.I(Mfifo_xin_raddr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3246 (
	.O(n3130),
	.I1(n3419),
	.I2(n2881), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3247 (
	.O(n3420),
	.I(Mfifo_xin_raddr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U3248 (
	.O(n3498),
	.I1(n3419),
	.I2(n3420),
	.I3(n3418), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3249 (
	.O(n3510),
	.I(n2882), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2X05AR9 U3250 (
	.O(n3131),
	.I1(n3498),
	.I2(n3510), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U3251 (
	.O(Mfifo_xin_M_rptr_rbinnext[3]),
	.B2(n3131),
	.I1(n3130), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3252 (
	.O(n3415),
	.I(Mfifo_coe_M_rptr_N1), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U3253 (
	.O(n3416),
	.B2(n3415),
	.I1(Mfifo_coe_raddr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3254 (
	.O(n2884),
	.I1(Mfifo_coe_raddr[1]),
	.I2(n3416), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3255 (
	.O(n3153),
	.I1(Mfifo_coe_raddr[1]),
	.I2(n3416), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U3256 (
	.O(Mfifo_coe_M_rptr_rbinnext[1]),
	.B2(n3153),
	.I1(n2884), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3257 (
	.O(n3325),
	.I(Mfifo_coe_raddr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3258 (
	.O(n3151),
	.I1(n3325),
	.I2(n2884), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA12X05AR9 U3259 (
	.O(Mfifo_coe_M_rptr_rbinnext[2]),
	.A1(n3151),
	.B1(n2884),
	.B2(n3325), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U3260 (
	.O(int_end_read),
	.I1(int_comp),
	.I2(n2883),
	.I3(n3101), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3261 (
	.O(n3324),
	.I(Mfifo_coe_raddr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3262 (
	.O(n3152),
	.A1(n3324),
	.B1(n3325),
	.B2(n2884), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3263 (
	.O(n3326),
	.I(Mfifo_coe_raddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U3264 (
	.O(n3406),
	.I1(n3326),
	.I2(n3324),
	.I3(n3325), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2X05AR9 U3265 (
	.O(n3150),
	.I1(n3406),
	.I2(n3416), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U3266 (
	.O(Mfifo_coe_M_rptr_rbinnext[3]),
	.B2(n3150),
	.I1(n3152), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3267 (
	.O(n3241),
	.I1(n2885),
	.I2(int_comp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3268 (
	.O(n3317),
	.I1(n3101),
	.I2(n3241), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3269 (
	.O(n3110),
	.I1(n3240),
	.I2(n3317), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3270 (
	.O(n3512),
	.A1(n3520),
	.B1(n2886),
	.B2(n3235), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3271 (
	.O(n2899),
	.I1(n3090),
	.I2(n3512), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3272 (
	.O(n2887),
	.I1(n2886),
	.I2(n3520), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3273 (
	.O(n3096),
	.A1(n2887),
	.B1(n3110),
	.B2(n2899), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3274 (
	.O(n3106),
	.I(n3110), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3275 (
	.O(n3129),
	.A1(n3106),
	.B1(n3091),
	.B2(n3096), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3276 (
	.O(n3126),
	.I(n3129), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3277 (
	.O(n3122),
	.I1(n2888),
	.I2(n2899), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3278 (
	.O(n2890),
	.I(n3122), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3279 (
	.O(n2889),
	.A1(n3119),
	.B1(Mcntl_Mcntldata_c_x_H[1]),
	.B2(Mcntl_Mcntldata_c_x_H[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3280 (
	.O(n2893),
	.A1(n3240),
	.B1(n3512),
	.B2(n2888), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3281 (
	.O(n2896),
	.I1(Mcntl_Mcntldata_x_H_reg[1]),
	.I2(Mcntl_Mcntldata_x_H_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3282 (
	.O(n2894),
	.A1(n2896),
	.B1(Mcntl_Mcntldata_x_H_reg[0]),
	.B2(Mcntl_Mcntldata_x_H_reg[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3283 (
	.O(n3113),
	.I(Mcntl_Mcntldata_x_H_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3284 (
	.O(n3112),
	.I1(n3113),
	.I2(n3087), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3285 (
	.O(n2897),
	.A1(n3317),
	.B1(n2888),
	.B2(n3090), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI222X05AR9 U3286 (
	.O(n2891),
	.A1(n2890),
	.A2(n2889),
	.B1(n2893),
	.B2(n2894),
	.C1(n3295),
	.C2(n2897), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA22X05AR9 U3287 (
	.O(n2085),
	.A1(n3126),
	.A2(Mcntl_Mcntldata_c_x_H[1]),
	.B1(n3129),
	.B2(n2891), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U3288 (
	.O(n2892),
	.I1(Mcntl_Mcntldata_x_H_reg[2]),
	.I2(Mcntl_Mcntldata_x_H_reg[1]),
	.I3(Mcntl_Mcntldata_x_H_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3289 (
	.O(n2898),
	.A1(n2892),
	.A2(Mcntl_Mcntldata_x_H_reg[3]),
	.B1B(n2892),
	.B2B(Mcntl_Mcntldata_x_H_reg[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3290 (
	.O(n3121),
	.I(n2893), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3291 (
	.O(n3117),
	.I(n2895), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3292 (
	.O(n3120),
	.A1(Mcntl_Mcntldata_x_H_reg[2]),
	.A2(n2896),
	.B1B(Mcntl_Mcntldata_x_H_reg[2]),
	.B2B(n2896), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3293 (
	.O(n3116),
	.I1(n3117),
	.I2(n3120), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3294 (
	.O(n3307),
	.A1(n3116),
	.A2(Mcntl_Mcntldata_x_H_reg[3]),
	.B1B(n3116),
	.B2B(n2898), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3295 (
	.O(n3125),
	.I(n2897), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3296 (
	.O(n2901),
	.A1(n2898),
	.A2(n3121),
	.B1(n3307),
	.B2(n3125), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3297 (
	.O(n3109),
	.I(n2899), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12B2X05AR9 U3298 (
	.O(n2900),
	.A1(n3126),
	.B1B(n3118),
	.B2B(n3109), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U3299 (
	.O(n2087),
	.A1(n3129),
	.A2(n2901),
	.B1B(Mcntl_Mcntldata_c_x_H[3]),
	.B2B(n2900), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3300 (
	.O(n3556),
	.I1(Mfifo_psum_waddr[2]),
	.I2(Mfifo_psum_waddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3301 (
	.O(n2904),
	.I1(n3547),
	.I2(Mfifo_psum_waddr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3302 (
	.O(n2902),
	.I1(n3547),
	.I2(Mfifo_psum_waddr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3303 (
	.O(Mfifo_psum_M_wptr_wbinnext[3]),
	.I1(n2904),
	.I2(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3304 (
	.O(n2903),
	.I1(Mfifo_psum_wptr[4]),
	.I2(n2902), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3305 (
	.O(Mfifo_psum_M_wptr_wbinnext[4]),
	.A1(n2903),
	.B1(Mfifo_psum_wptr[4]),
	.B2(n2902), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA22X05AR9 U3306 (
	.O(Mfifo_psum_M_wptr_wgraynext[3]),
	.A1(Mfifo_psum_M_wptr_wbinnext[3]),
	.A2(Mfifo_psum_M_wptr_wbinnext[4]),
	.B1(n2904),
	.B2(n2903), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3307 (
	.O(n3316),
	.I1(Mcntl_Mcntldata_c_p_wd4[0]),
	.I2(n3839), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3308 (
	.O(n3315),
	.I(Mcntl_Mcntldata_c_p_wd4[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3309 (
	.O(n3311),
	.I1(n3316),
	.I2(n3315), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U3310 (
	.O(n3319),
	.B2(n3311),
	.I1(n3181), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3311 (
	.O(n3280),
	.I1(n2905),
	.I2(int_send), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3312 (
	.O(n3263),
	.I(n3280), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3313 (
	.O(n3183),
	.I1(n3319),
	.I2(n3263), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2X05AR9 U3314 (
	.O(n2906),
	.I1(n3183),
	.I2(n2907), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3315 (
	.O(n2925),
	.I1(n3147),
	.I2(n2906), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2B1X05AR9 U3316 (
	.O(n2908),
	.B2(n3183),
	.I1(n2907), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3317 (
	.O(n2923),
	.I1(n2908),
	.I2(n3147), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U3318 (
	.O(n2077),
	.A1(n2925),
	.A2(n2909),
	.B1B(C175_DATA2_0),
	.B2B(n2923), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3319 (
	.O(n2910),
	.I(DP_OP_1207J5_130_8771_n6), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U3320 (
	.O(n2076),
	.A1(n2925),
	.A2(n2913),
	.B1B(C175_DATA2_2),
	.B2B(n2923), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3321 (
	.O(n2918),
	.I(x_addr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3322 (
	.O(n2916),
	.I1(n2915),
	.I2(n2914), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3323 (
	.O(n2917),
	.I(n2916), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3324 (
	.O(n3205),
	.I1(n2917),
	.I2(n3110), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U3325 (
	.O(n2071),
	.A1(n2918),
	.A2(n3205),
	.B1B(C174_DATA2_0),
	.B2B(n2916), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U3326 (
	.O(n2075),
	.A1(n2925),
	.A2(n3209),
	.B1B(C175_DATA2_3),
	.B2B(n2923), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3327 (
	.O(n2919),
	.I(x_addr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U3328 (
	.O(n2074),
	.A1(n2925),
	.A2(n2920),
	.B1B(C175_DATA2_4),
	.B2B(n2923), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3329 (
	.O(n2921),
	.I(x_addr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U3330 (
	.O(n2070),
	.A1(n2921),
	.A2(n3205),
	.B1B(C174_DATA2_2),
	.B2B(n2916), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   XOR2X05AR9 U3331 (
	.O(n2922),
	.I1(n3843),
	.I2(Mcntl_Mcntldata_N453), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   XOR2X05AR9 U3332 (
	.O(n2924),
	.I1(DP_OP_1207J5_130_8771_n2),
	.I2(n2922), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U3333 (
	.O(n2073),
	.A1(n3208),
	.A2(n2925),
	.B1B(n2924),
	.B2B(n2923), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2X05AR9 U3334 (
	.O(n3833),
	.I1(psum_addr[1]),
	.I2(DP_OP_1207J5_130_8771_n6), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3335 (
	.O(n2926),
	.I(x_addr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U3336 (
	.O(n2069),
	.A1(n2926),
	.A2(n3205),
	.B1B(C174_DATA2_3),
	.B2B(n2916), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3337 (
	.O(n2927),
	.I(x_addr[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U3338 (
	.O(n2068),
	.A1(n2927),
	.A2(n3205),
	.B1B(C174_DATA2_4),
	.B2B(n2916), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3339 (
	.O(n2928),
	.I(x_addr[5]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22B2X05AR9 U3340 (
	.O(n2067),
	.A1(n2928),
	.A2(n3205),
	.B1B(C174_DATA2_5),
	.B2B(n2916), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3341 (
	.O(n3523),
	.I(Mcntl_Mcntldata_x_W_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3342 (
	.O(n3514),
	.I(Mcntl_Mcntldata_x_W_reg[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3343 (
	.O(n3513),
	.I1(n3523),
	.I2(n3514), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2X05AR9 U3344 (
	.O(n2930),
	.I1(n3513),
	.I2(Mcntl_Mcntldata_x_W_reg[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3345 (
	.O(n3186),
	.I(Mcntl_Mcntldata_x_W_reg[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3346 (
	.O(n2929),
	.I1(n3513),
	.I2(n3186), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3347 (
	.O(n3093),
	.I1(n2930),
	.I2(n2929), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3348 (
	.O(n3310),
	.I1(n3513),
	.I2(Mcntl_Mcntldata_x_W_reg[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3349 (
	.O(n3258),
	.I(Mcntl_Mcntldata_x_W_reg[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3350 (
	.O(n2931),
	.I1(n3310),
	.I2(n3258), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3351 (
	.O(n3312),
	.A1(n2931),
	.B1(n3093),
	.B2(n3310), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3352 (
	.O(n2961),
	.I1(n3310),
	.I2(Mcntl_Mcntldata_ky_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3353 (
	.O(n2938),
	.I(n2961), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U3354 (
	.O(n2950),
	.I1(n3312),
	.I2(Mcntl_Mcntldata_ky_reg[1]),
	.I3(n2938), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3355 (
	.O(n2932),
	.I(n3310), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U3356 (
	.O(n2933),
	.I1(n2932),
	.I2(Mcntl_Mcntldata_ky_reg[1]),
	.I3(Mcntl_Mcntldata_x_W_reg[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3357 (
	.O(n2939),
	.I1(n2950),
	.I2(n2933), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3358 (
	.O(n2935),
	.I1(n3312),
	.I2(Mcntl_Mcntldata_ky_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3359 (
	.O(n2934),
	.I1(n3310),
	.I2(Mcntl_Mcntldata_ky_reg[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3360 (
	.O(n2951),
	.I1(n2935),
	.I2(n2934), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3361 (
	.O(n2937),
	.I1(n3312),
	.I2(Mcntl_Mcntldata_ky_reg[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3362 (
	.O(n2936),
	.I1(Mcntl_Mcntldata_ky_reg[0]),
	.I2(Mcntl_Mcntldata_x_W_reg[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3363 (
	.O(n2943),
	.I1(n2937),
	.I2(n2936), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U3364 (
	.O(n2944),
	.I1(n2951),
	.I2(n2943),
	.I3(n2938), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   XNOR2X05AR9 U3365 (
	.O(n2941),
	.I1(n2939),
	.I2(n2944), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3366 (
	.O(n2940),
	.I(n2939), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3367 (
	.O(n2942),
	.A1(n2941),
	.A2(n2947),
	.B1(n2959),
	.B2(n2940), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   XOR2X05AR9 U3368 (
	.O(DP_OP_1205J5_125_5849_n12),
	.I1(n2942),
	.I2(C2_Z_0), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3369 (
	.O(n2948),
	.I1(n2943),
	.I2(n2961), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3370 (
	.O(n2945),
	.I(n2948), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3371 (
	.O(n2946),
	.A1(n2944),
	.B1(n2945),
	.B2(n2951), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3372 (
	.O(n2949),
	.A1(n2959),
	.A2(n2948),
	.B1(n2947),
	.B2(n2946), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   XOR2X05AR9 U3373 (
	.O(DP_OP_1205J5_125_5849_n13),
	.I1(n2949),
	.I2(C2_Z_0), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3374 (
	.O(n2956),
	.I1(n2951),
	.I2(n2950), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   MUX2BX05AR9 U3375 (
	.OB(n2954),
	.I0(n2956),
	.I1(n2951),
	.S(n2961), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3376 (
	.O(n2952),
	.I(n3165), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3377 (
	.O(n3313),
	.I(n3093), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3378 (
	.O(n2955),
	.A1(n2954),
	.A2(n2962),
	.B1(n2958),
	.B2(n3313), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3379 (
	.O(n2957),
	.A1(n2955),
	.B1(n2959),
	.B2(n2956), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3380 (
	.O(n2965),
	.I(n2958), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3381 (
	.O(n2964),
	.A1(n2960),
	.B1(n2962),
	.B2(n2961), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3382 (
	.O(n2966),
	.A1(n2964),
	.B1(n2963),
	.C1(n2965),
	.C2(n3310), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3383 (
	.O(n3048),
	.I1(Mfifo_xin_waddr[1]),
	.I2(Mfifo_xin_waddr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3384 (
	.O(n2973),
	.I(Mfifo_xin_waddr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3385 (
	.O(n3005),
	.I(ext_xin[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3386 (
	.O(n2213),
	.A1(n2967),
	.A2(n3005),
	.B1B(n2967),
	.B2B(Mfifo_xin_M_ffmem_mem_14__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3387 (
	.O(n3001),
	.I(ext_xin[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3388 (
	.O(n2211),
	.A1(n2967),
	.A2(n3001),
	.B1B(n2967),
	.B2B(Mfifo_xin_M_ffmem_mem_14__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3389 (
	.O(n3004),
	.I(ext_xin[5]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3390 (
	.O(n2214),
	.A1(n2967),
	.A2(n3004),
	.B1B(n2967),
	.B2B(Mfifo_xin_M_ffmem_mem_14__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3391 (
	.O(n3002),
	.I(ext_xin[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3392 (
	.O(n2210),
	.A1(n2967),
	.A2(n3002),
	.B1B(n2967),
	.B2B(Mfifo_xin_M_ffmem_mem_14__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3393 (
	.O(n2999),
	.I(ext_xin[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3394 (
	.O(n2215),
	.A1(n2967),
	.A2(n2999),
	.B1B(n2967),
	.B2B(Mfifo_xin_M_ffmem_mem_14__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3395 (
	.O(n3003),
	.I(ext_xin[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3396 (
	.O(n2212),
	.A1(n2967),
	.A2(n3003),
	.B1B(n2967),
	.B2B(Mfifo_xin_M_ffmem_mem_14__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3397 (
	.O(n2997),
	.I(ext_xin[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3398 (
	.O(n2217),
	.A1(n2967),
	.A2(n2997),
	.B1B(n2967),
	.B2B(Mfifo_xin_M_ffmem_mem_14__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3399 (
	.O(n2998),
	.I(ext_xin[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3400 (
	.O(n2216),
	.A1(n2967),
	.A2(n2998),
	.B1B(n2967),
	.B2B(Mfifo_xin_M_ffmem_mem_14__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3401 (
	.O(n3066),
	.I1(Mfifo_coe_waddr[1]),
	.I2(Mfifo_coe_waddr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3402 (
	.O(n3019),
	.I(ext_coe[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3403 (
	.O(n2292),
	.A1(n3067),
	.A2(n3019),
	.B1B(Mfifo_coe_M_ffmem_mem_7__3_),
	.B2B(n3067), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3404 (
	.O(n3023),
	.I(ext_coe[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3405 (
	.O(n2290),
	.A1(n3067),
	.A2(n3023),
	.B1B(Mfifo_coe_M_ffmem_mem_7__1_),
	.B2B(n3067), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3406 (
	.O(n2295),
	.A1(n3067),
	.A2(n3027),
	.B1B(Mfifo_coe_M_ffmem_mem_7__6_),
	.B2B(n3067), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3407 (
	.O(n3026),
	.I(ext_coe[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3408 (
	.O(n2293),
	.A1(n3067),
	.A2(n3026),
	.B1B(Mfifo_coe_M_ffmem_mem_7__4_),
	.B2B(n3067), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3409 (
	.O(n3020),
	.I(ext_coe[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3410 (
	.O(n2296),
	.A1(n3067),
	.A2(n3020),
	.B1B(Mfifo_coe_M_ffmem_mem_7__7_),
	.B2B(n3067), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3411 (
	.O(n3025),
	.I(ext_coe[5]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3412 (
	.O(n2294),
	.A1(n3067),
	.A2(n3025),
	.B1B(Mfifo_coe_M_ffmem_mem_7__5_),
	.B2B(n3067), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3413 (
	.O(n3017),
	.I(ext_coe[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3414 (
	.O(n2297),
	.A1(n3067),
	.A2(n3017),
	.B1B(Mfifo_coe_M_ffmem_mem_7__0_),
	.B2B(n3067), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3415 (
	.O(n3021),
	.I(ext_coe[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3416 (
	.O(n2291),
	.A1(n3067),
	.A2(n3021),
	.B1B(Mfifo_coe_M_ffmem_mem_7__2_),
	.B2B(n3067), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3417 (
	.O(n2994),
	.I1(Mfifo_xin_waddr[2]),
	.I2(n3055), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U3418 (
	.O(n2972),
	.I1(n2969),
	.I2(n2994), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3419 (
	.O(n2199),
	.A1(n2972),
	.A2(n2999),
	.B1B(n2972),
	.B2B(Mfifo_xin_M_ffmem_mem_12__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3420 (
	.O(n2198),
	.A1(n2972),
	.A2(n3004),
	.B1B(n2972),
	.B2B(Mfifo_xin_M_ffmem_mem_12__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3421 (
	.O(n2968),
	.I(Mfifo_xin_waddr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3422 (
	.O(n2993),
	.I1(n3055),
	.I2(n2968), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U3423 (
	.O(n2971),
	.I1(n2969),
	.I2(n2993), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3424 (
	.O(n2163),
	.A1(n2971),
	.A2(n3001),
	.B1B(n2971),
	.B2B(Mfifo_xin_M_ffmem_mem_8__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3425 (
	.O(n2200),
	.A1(n2972),
	.A2(n2998),
	.B1B(n2972),
	.B2B(Mfifo_xin_M_ffmem_mem_12__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3426 (
	.O(n2165),
	.A1(n2971),
	.A2(n3005),
	.B1B(n2971),
	.B2B(Mfifo_xin_M_ffmem_mem_8__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3427 (
	.O(n2166),
	.A1(n2971),
	.A2(n3004),
	.B1B(n2971),
	.B2B(Mfifo_xin_M_ffmem_mem_8__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3428 (
	.O(n2167),
	.A1(n2971),
	.A2(n2999),
	.B1B(n2971),
	.B2B(Mfifo_xin_M_ffmem_mem_8__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3429 (
	.O(n2168),
	.A1(n2971),
	.A2(n2998),
	.B1B(n2971),
	.B2B(Mfifo_xin_M_ffmem_mem_8__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3430 (
	.O(n2169),
	.A1(n2971),
	.A2(n2997),
	.B1B(n2971),
	.B2B(Mfifo_xin_M_ffmem_mem_8__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3431 (
	.O(n2992),
	.I1(Mfifo_xin_waddr[1]),
	.I2(n2968), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U3432 (
	.O(n2970),
	.I1(n2969),
	.I2(n2992), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3433 (
	.O(n2178),
	.A1(n2970),
	.A2(n3002),
	.B1B(n2970),
	.B2B(Mfifo_xin_M_ffmem_mem_10__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3434 (
	.O(n2179),
	.A1(n2970),
	.A2(n3001),
	.B1B(n2970),
	.B2B(Mfifo_xin_M_ffmem_mem_10__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3435 (
	.O(n2180),
	.A1(n2970),
	.A2(n3003),
	.B1B(n2970),
	.B2B(Mfifo_xin_M_ffmem_mem_10__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3436 (
	.O(n2181),
	.A1(n2970),
	.A2(n3005),
	.B1B(n2970),
	.B2B(Mfifo_xin_M_ffmem_mem_10__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3437 (
	.O(n2197),
	.A1(n2972),
	.A2(n3005),
	.B1B(n2972),
	.B2B(Mfifo_xin_M_ffmem_mem_12__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3438 (
	.O(n2182),
	.A1(n2970),
	.A2(n3004),
	.B1B(n2970),
	.B2B(Mfifo_xin_M_ffmem_mem_10__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3439 (
	.O(n2185),
	.A1(n2970),
	.A2(n2997),
	.B1B(n2970),
	.B2B(Mfifo_xin_M_ffmem_mem_10__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3440 (
	.O(n2183),
	.A1(n2970),
	.A2(n2999),
	.B1B(n2970),
	.B2B(Mfifo_xin_M_ffmem_mem_10__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3441 (
	.O(n2201),
	.A1(n2972),
	.A2(n2997),
	.B1B(n2972),
	.B2B(Mfifo_xin_M_ffmem_mem_12__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3442 (
	.O(n2184),
	.A1(n2970),
	.A2(n2998),
	.B1B(n2970),
	.B2B(Mfifo_xin_M_ffmem_mem_10__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3443 (
	.O(n2164),
	.A1(n2971),
	.A2(n3003),
	.B1B(n2971),
	.B2B(Mfifo_xin_M_ffmem_mem_8__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3444 (
	.O(n2194),
	.A1(n2972),
	.A2(n3002),
	.B1B(n2972),
	.B2B(Mfifo_xin_M_ffmem_mem_12__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3445 (
	.O(n2162),
	.A1(n2971),
	.A2(n3002),
	.B1B(n2971),
	.B2B(Mfifo_xin_M_ffmem_mem_8__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3446 (
	.O(n2195),
	.A1(n2972),
	.A2(n3001),
	.B1B(n2972),
	.B2B(Mfifo_xin_M_ffmem_mem_12__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3447 (
	.O(n2196),
	.A1(n2972),
	.A2(n3003),
	.B1B(n2972),
	.B2B(Mfifo_xin_M_ffmem_mem_12__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X1AR9 U3448 (
	.O(n2985),
	.I1(Mfifo_coe_waddr[3]),
	.I2(n3222), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3449 (
	.O(n2359),
	.A1(n3064),
	.A2(n3027),
	.B1B(Mfifo_coe_M_ffmem_mem_15__6_),
	.B2B(n3064), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3450 (
	.O(n2357),
	.A1(n3064),
	.A2(n3026),
	.B1B(Mfifo_coe_M_ffmem_mem_15__4_),
	.B2B(n3064), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3451 (
	.O(n2360),
	.A1(n3064),
	.A2(n3020),
	.B1B(Mfifo_coe_M_ffmem_mem_15__7_),
	.B2B(n3064), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3452 (
	.O(n2358),
	.A1(n3064),
	.A2(n3025),
	.B1B(Mfifo_coe_M_ffmem_mem_15__5_),
	.B2B(n3064), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3453 (
	.O(n2355),
	.A1(n3064),
	.A2(n3021),
	.B1B(Mfifo_coe_M_ffmem_mem_15__2_),
	.B2B(n3064), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3454 (
	.O(n2354),
	.A1(n3064),
	.A2(n3023),
	.B1B(Mfifo_coe_M_ffmem_mem_15__1_),
	.B2B(n3064), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3455 (
	.O(n2356),
	.A1(n3064),
	.A2(n3019),
	.B1B(Mfifo_coe_M_ffmem_mem_15__3_),
	.B2B(n3064), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3456 (
	.O(n2361),
	.A1(n3064),
	.A2(n3017),
	.B1B(Mfifo_coe_M_ffmem_mem_15__0_),
	.B2B(n3064), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3457 (
	.O(n2120),
	.A1(n2977),
	.A2(n2998),
	.B1B(n2977),
	.B2B(Mfifo_xin_M_ffmem_mem_2__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3458 (
	.O(n2103),
	.A1(n2974),
	.A2(n2999),
	.B1B(n2974),
	.B2B(Mfifo_xin_M_ffmem_mem_0__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3459 (
	.O(n2101),
	.A1(n2974),
	.A2(n3005),
	.B1B(n2974),
	.B2B(Mfifo_xin_M_ffmem_mem_0__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3460 (
	.O(n2102),
	.A1(n2974),
	.A2(n3004),
	.B1B(n2974),
	.B2B(Mfifo_xin_M_ffmem_mem_0__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3461 (
	.O(n2116),
	.A1(n2977),
	.A2(n3003),
	.B1B(n2977),
	.B2B(Mfifo_xin_M_ffmem_mem_2__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3462 (
	.O(n2104),
	.A1(n2974),
	.A2(n2998),
	.B1B(n2974),
	.B2B(Mfifo_xin_M_ffmem_mem_0__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3463 (
	.O(n2132),
	.A1(n2975),
	.A2(n3003),
	.B1B(n2975),
	.B2B(Mfifo_xin_M_ffmem_mem_4__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3464 (
	.O(n2114),
	.A1(n2977),
	.A2(n3002),
	.B1B(n2977),
	.B2B(Mfifo_xin_M_ffmem_mem_2__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3465 (
	.O(n2135),
	.A1(n2975),
	.A2(n2999),
	.B1B(n2975),
	.B2B(Mfifo_xin_M_ffmem_mem_4__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3466 (
	.O(n2121),
	.A1(n2977),
	.A2(n2997),
	.B1B(n2977),
	.B2B(Mfifo_xin_M_ffmem_mem_2__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3467 (
	.O(n2130),
	.A1(n2975),
	.A2(n3002),
	.B1B(n2975),
	.B2B(Mfifo_xin_M_ffmem_mem_4__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3468 (
	.O(n2105),
	.A1(n2974),
	.A2(n2997),
	.B1B(n2974),
	.B2B(Mfifo_xin_M_ffmem_mem_0__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3469 (
	.O(n2136),
	.A1(n2975),
	.A2(n2998),
	.B1B(n2975),
	.B2B(Mfifo_xin_M_ffmem_mem_4__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3470 (
	.O(n2133),
	.A1(n2975),
	.A2(n3005),
	.B1B(n2975),
	.B2B(Mfifo_xin_M_ffmem_mem_4__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3471 (
	.O(n2115),
	.A1(n2977),
	.A2(n3001),
	.B1B(n2977),
	.B2B(Mfifo_xin_M_ffmem_mem_2__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3472 (
	.O(n2134),
	.A1(n2975),
	.A2(n3004),
	.B1B(n2975),
	.B2B(Mfifo_xin_M_ffmem_mem_4__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3473 (
	.O(n2131),
	.A1(n2975),
	.A2(n3001),
	.B1B(n2975),
	.B2B(Mfifo_xin_M_ffmem_mem_4__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3474 (
	.O(n2118),
	.A1(n2977),
	.A2(n3004),
	.B1B(n2977),
	.B2B(Mfifo_xin_M_ffmem_mem_2__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3475 (
	.O(n2119),
	.A1(n2977),
	.A2(n2999),
	.B1B(n2977),
	.B2B(Mfifo_xin_M_ffmem_mem_2__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3476 (
	.O(n2098),
	.A1(n2974),
	.A2(n3002),
	.B1B(n2974),
	.B2B(Mfifo_xin_M_ffmem_mem_0__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3477 (
	.O(n2099),
	.A1(n2974),
	.A2(n3001),
	.B1B(n2974),
	.B2B(Mfifo_xin_M_ffmem_mem_0__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3478 (
	.O(n2100),
	.A1(n2974),
	.A2(n3003),
	.B1B(n2974),
	.B2B(Mfifo_xin_M_ffmem_mem_0__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3479 (
	.O(n2137),
	.A1(n2975),
	.A2(n2997),
	.B1B(n2975),
	.B2B(Mfifo_xin_M_ffmem_mem_4__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3480 (
	.O(n2146),
	.A1(n2978),
	.A2(n3002),
	.B1B(n2978),
	.B2B(Mfifo_xin_M_ffmem_mem_6__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3481 (
	.O(n2147),
	.A1(n2978),
	.A2(n3001),
	.B1B(n2978),
	.B2B(Mfifo_xin_M_ffmem_mem_6__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3482 (
	.O(n2148),
	.A1(n2978),
	.A2(n3003),
	.B1B(n2978),
	.B2B(Mfifo_xin_M_ffmem_mem_6__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3483 (
	.O(n2117),
	.A1(n2977),
	.A2(n3005),
	.B1B(n2977),
	.B2B(Mfifo_xin_M_ffmem_mem_2__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3484 (
	.O(n2149),
	.A1(n2978),
	.A2(n3005),
	.B1B(n2978),
	.B2B(Mfifo_xin_M_ffmem_mem_6__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3485 (
	.O(n2150),
	.A1(n2978),
	.A2(n3004),
	.B1B(n2978),
	.B2B(Mfifo_xin_M_ffmem_mem_6__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3486 (
	.O(n2151),
	.A1(n2978),
	.A2(n2999),
	.B1B(n2978),
	.B2B(Mfifo_xin_M_ffmem_mem_6__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3487 (
	.O(n2152),
	.A1(n2978),
	.A2(n2998),
	.B1B(n2978),
	.B2B(Mfifo_xin_M_ffmem_mem_6__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3488 (
	.O(n2153),
	.A1(n2978),
	.A2(n2997),
	.B1B(n2978),
	.B2B(Mfifo_xin_M_ffmem_mem_6__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3489 (
	.O(n3014),
	.I1(Mfifo_coe_waddr[2]),
	.I2(n3071), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U3490 (
	.O(n2983),
	.I1(n2981),
	.I2(n3014), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3491 (
	.O(n2281),
	.A1(n2983),
	.A2(n3017),
	.B1B(n2983),
	.B2B(Mfifo_coe_M_ffmem_mem_5__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3492 (
	.O(n2280),
	.A1(n2983),
	.A2(n3020),
	.B1B(n2983),
	.B2B(Mfifo_coe_M_ffmem_mem_5__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3493 (
	.O(n2279),
	.A1(n2983),
	.A2(n3027),
	.B1B(n2983),
	.B2B(Mfifo_coe_M_ffmem_mem_5__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U3494 (
	.O(n2986),
	.I1(n2985),
	.I2(n3014), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3495 (
	.O(n2345),
	.A1(n2986),
	.A2(n3017),
	.B1B(n2986),
	.B2B(Mfifo_coe_M_ffmem_mem_13__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3496 (
	.O(n2277),
	.A1(n2983),
	.A2(n3026),
	.B1B(n2983),
	.B2B(Mfifo_coe_M_ffmem_mem_5__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3497 (
	.O(n2276),
	.A1(n2983),
	.A2(n3019),
	.B1B(n2983),
	.B2B(Mfifo_coe_M_ffmem_mem_5__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3498 (
	.O(n2275),
	.A1(n2983),
	.A2(n3021),
	.B1B(n2983),
	.B2B(Mfifo_coe_M_ffmem_mem_5__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3499 (
	.O(n2274),
	.A1(n2983),
	.A2(n3023),
	.B1B(n2983),
	.B2B(Mfifo_coe_M_ffmem_mem_5__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3500 (
	.O(n2980),
	.I(Mfifo_coe_waddr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3501 (
	.O(n3016),
	.I1(Mfifo_coe_waddr[1]),
	.I2(n2980), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U3502 (
	.O(n2979),
	.I1(n2981),
	.I2(n3016), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3503 (
	.O(n2265),
	.A1(n2979),
	.A2(n3017),
	.B1B(n2979),
	.B2B(Mfifo_coe_M_ffmem_mem_3__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3504 (
	.O(n2264),
	.A1(n2979),
	.A2(n3020),
	.B1B(n2979),
	.B2B(Mfifo_coe_M_ffmem_mem_3__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3505 (
	.O(n2263),
	.A1(n2979),
	.A2(n3027),
	.B1B(n2979),
	.B2B(Mfifo_coe_M_ffmem_mem_3__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3506 (
	.O(n2262),
	.A1(n2979),
	.A2(n3025),
	.B1B(n2979),
	.B2B(Mfifo_coe_M_ffmem_mem_3__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3507 (
	.O(n2261),
	.A1(n2979),
	.A2(n3026),
	.B1B(n2979),
	.B2B(Mfifo_coe_M_ffmem_mem_3__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3508 (
	.O(n2260),
	.A1(n2979),
	.A2(n3019),
	.B1B(n2979),
	.B2B(Mfifo_coe_M_ffmem_mem_3__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3509 (
	.O(n2259),
	.A1(n2979),
	.A2(n3021),
	.B1B(n2979),
	.B2B(Mfifo_coe_M_ffmem_mem_3__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3510 (
	.O(n2258),
	.A1(n2979),
	.A2(n3023),
	.B1B(n2979),
	.B2B(Mfifo_coe_M_ffmem_mem_3__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3511 (
	.O(n2344),
	.A1(n2986),
	.A2(n3020),
	.B1B(n2986),
	.B2B(Mfifo_coe_M_ffmem_mem_13__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3512 (
	.O(n3013),
	.I1(n3071),
	.I2(n2980), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3513 (
	.O(n2249),
	.A1(n2982),
	.A2(n3017),
	.B1B(n2982),
	.B2B(Mfifo_coe_M_ffmem_mem_1__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3514 (
	.O(n2248),
	.A1(n2982),
	.A2(n3020),
	.B1B(n2982),
	.B2B(Mfifo_coe_M_ffmem_mem_1__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3515 (
	.O(n2343),
	.A1(n2986),
	.A2(n3027),
	.B1B(n2986),
	.B2B(Mfifo_coe_M_ffmem_mem_13__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3516 (
	.O(n2247),
	.A1(n2982),
	.A2(n3027),
	.B1B(n2982),
	.B2B(Mfifo_coe_M_ffmem_mem_1__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3517 (
	.O(n2246),
	.A1(n2982),
	.A2(n3025),
	.B1B(n2982),
	.B2B(Mfifo_coe_M_ffmem_mem_1__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3518 (
	.O(n2245),
	.A1(n2982),
	.A2(n3026),
	.B1B(n2982),
	.B2B(Mfifo_coe_M_ffmem_mem_1__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3519 (
	.O(n2244),
	.A1(n2982),
	.A2(n3019),
	.B1B(n2982),
	.B2B(Mfifo_coe_M_ffmem_mem_1__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3520 (
	.O(n2243),
	.A1(n2982),
	.A2(n3021),
	.B1B(n2982),
	.B2B(Mfifo_coe_M_ffmem_mem_1__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3521 (
	.O(n2242),
	.A1(n2982),
	.A2(n3023),
	.B1B(n2982),
	.B2B(Mfifo_coe_M_ffmem_mem_1__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3522 (
	.O(n2342),
	.A1(n2986),
	.A2(n3025),
	.B1B(n2986),
	.B2B(Mfifo_coe_M_ffmem_mem_13__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3523 (
	.O(n2278),
	.A1(n2983),
	.A2(n3025),
	.B1B(n2983),
	.B2B(Mfifo_coe_M_ffmem_mem_5__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3524 (
	.O(n2341),
	.A1(n2986),
	.A2(n3026),
	.B1B(n2986),
	.B2B(Mfifo_coe_M_ffmem_mem_13__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3525 (
	.O(n2340),
	.A1(n2986),
	.A2(n3019),
	.B1B(n2986),
	.B2B(Mfifo_coe_M_ffmem_mem_13__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U3526 (
	.O(n2984),
	.I1(n2985),
	.I2(n3013), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3527 (
	.O(n2306),
	.A1(n2984),
	.A2(n3023),
	.B1B(n2984),
	.B2B(Mfifo_coe_M_ffmem_mem_9__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3528 (
	.O(n2307),
	.A1(n2984),
	.A2(n3021),
	.B1B(n2984),
	.B2B(Mfifo_coe_M_ffmem_mem_9__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3529 (
	.O(n2308),
	.A1(n2984),
	.A2(n3019),
	.B1B(n2984),
	.B2B(Mfifo_coe_M_ffmem_mem_9__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3530 (
	.O(n2309),
	.A1(n2984),
	.A2(n3026),
	.B1B(n2984),
	.B2B(Mfifo_coe_M_ffmem_mem_9__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3531 (
	.O(n2310),
	.A1(n2984),
	.A2(n3025),
	.B1B(n2984),
	.B2B(Mfifo_coe_M_ffmem_mem_9__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3532 (
	.O(n2311),
	.A1(n2984),
	.A2(n3027),
	.B1B(n2984),
	.B2B(Mfifo_coe_M_ffmem_mem_9__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3533 (
	.O(n2312),
	.A1(n2984),
	.A2(n3020),
	.B1B(n2984),
	.B2B(Mfifo_coe_M_ffmem_mem_9__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3534 (
	.O(n2313),
	.A1(n2984),
	.A2(n3017),
	.B1B(n2984),
	.B2B(Mfifo_coe_M_ffmem_mem_9__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U3535 (
	.O(n2987),
	.I1(n2985),
	.I2(n3016), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3536 (
	.O(n2322),
	.A1(n2987),
	.A2(n3023),
	.B1B(n2987),
	.B2B(Mfifo_coe_M_ffmem_mem_11__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3537 (
	.O(n2323),
	.A1(n2987),
	.A2(n3021),
	.B1B(n2987),
	.B2B(Mfifo_coe_M_ffmem_mem_11__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3538 (
	.O(n2324),
	.A1(n2987),
	.A2(n3019),
	.B1B(n2987),
	.B2B(Mfifo_coe_M_ffmem_mem_11__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3539 (
	.O(n2325),
	.A1(n2987),
	.A2(n3026),
	.B1B(n2987),
	.B2B(Mfifo_coe_M_ffmem_mem_11__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3540 (
	.O(n2339),
	.A1(n2986),
	.A2(n3021),
	.B1B(n2986),
	.B2B(Mfifo_coe_M_ffmem_mem_13__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3541 (
	.O(n2327),
	.A1(n2987),
	.A2(n3027),
	.B1B(n2987),
	.B2B(Mfifo_coe_M_ffmem_mem_11__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3542 (
	.O(n2328),
	.A1(n2987),
	.A2(n3020),
	.B1B(n2987),
	.B2B(Mfifo_coe_M_ffmem_mem_11__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3543 (
	.O(n2329),
	.A1(n2987),
	.A2(n3017),
	.B1B(n2987),
	.B2B(Mfifo_coe_M_ffmem_mem_11__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3544 (
	.O(n2338),
	.A1(n2986),
	.A2(n3023),
	.B1B(n2986),
	.B2B(Mfifo_coe_M_ffmem_mem_13__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3545 (
	.O(n2326),
	.A1(n2987),
	.A2(n3025),
	.B1B(n2987),
	.B2B(Mfifo_coe_M_ffmem_mem_11__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3546 (
	.O(n2154),
	.A1(n3050),
	.A2(n3002),
	.B1B(Mfifo_xin_M_ffmem_mem_7__1_),
	.B2B(n3050), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3547 (
	.O(n2155),
	.A1(n3050),
	.A2(n3001),
	.B1B(Mfifo_xin_M_ffmem_mem_7__2_),
	.B2B(n3050), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3548 (
	.O(n2156),
	.A1(n3050),
	.A2(n3003),
	.B1B(Mfifo_xin_M_ffmem_mem_7__3_),
	.B2B(n3050), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3549 (
	.O(n2157),
	.A1(n3050),
	.A2(n3005),
	.B1B(Mfifo_xin_M_ffmem_mem_7__4_),
	.B2B(n3050), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3550 (
	.O(n2158),
	.A1(n3050),
	.A2(n3004),
	.B1B(Mfifo_xin_M_ffmem_mem_7__5_),
	.B2B(n3050), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3551 (
	.O(n2159),
	.A1(n3050),
	.A2(n2999),
	.B1B(Mfifo_xin_M_ffmem_mem_7__6_),
	.B2B(n3050), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3552 (
	.O(n2160),
	.A1(n3050),
	.A2(n2998),
	.B1B(Mfifo_xin_M_ffmem_mem_7__7_),
	.B2B(n3050), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3553 (
	.O(n2161),
	.A1(n3050),
	.A2(n2997),
	.B1B(Mfifo_xin_M_ffmem_mem_7__0_),
	.B2B(n3050), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X1AR9 U3554 (
	.O(n2989),
	.I1(Mfifo_xin_waddr[3]),
	.I2(n3213), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3555 (
	.O(n2223),
	.A1(n3051),
	.A2(n2999),
	.B1B(Mfifo_xin_M_ffmem_mem_15__6_),
	.B2B(n3051), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3556 (
	.O(n2219),
	.A1(n3051),
	.A2(n3001),
	.B1B(Mfifo_xin_M_ffmem_mem_15__2_),
	.B2B(n3051), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3557 (
	.O(n2225),
	.A1(n3051),
	.A2(n2997),
	.B1B(Mfifo_xin_M_ffmem_mem_15__0_),
	.B2B(n3051), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3558 (
	.O(n2224),
	.A1(n3051),
	.A2(n2998),
	.B1B(Mfifo_xin_M_ffmem_mem_15__7_),
	.B2B(n3051), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3559 (
	.O(n2220),
	.A1(n3051),
	.A2(n3003),
	.B1B(Mfifo_xin_M_ffmem_mem_15__3_),
	.B2B(n3051), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3560 (
	.O(n2222),
	.A1(n3051),
	.A2(n3004),
	.B1B(Mfifo_xin_M_ffmem_mem_15__5_),
	.B2B(n3051), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3561 (
	.O(n2221),
	.A1(n3051),
	.A2(n3005),
	.B1B(Mfifo_xin_M_ffmem_mem_15__4_),
	.B2B(n3051), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3562 (
	.O(n2218),
	.A1(n3051),
	.A2(n3002),
	.B1B(Mfifo_xin_M_ffmem_mem_15__1_),
	.B2B(n3051), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3563 (
	.O(n2171),
	.A1(n2988),
	.A2(n3001),
	.B1B(n2988),
	.B2B(Mfifo_xin_M_ffmem_mem_9__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3564 (
	.O(n2172),
	.A1(n2988),
	.A2(n3003),
	.B1B(n2988),
	.B2B(Mfifo_xin_M_ffmem_mem_9__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3565 (
	.O(n2170),
	.A1(n2988),
	.A2(n3002),
	.B1B(n2988),
	.B2B(Mfifo_xin_M_ffmem_mem_9__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3566 (
	.O(n2174),
	.A1(n2988),
	.A2(n3004),
	.B1B(n2988),
	.B2B(Mfifo_xin_M_ffmem_mem_9__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3567 (
	.O(n2175),
	.A1(n2988),
	.A2(n2999),
	.B1B(n2988),
	.B2B(Mfifo_xin_M_ffmem_mem_9__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3568 (
	.O(n2173),
	.A1(n2988),
	.A2(n3005),
	.B1B(n2988),
	.B2B(Mfifo_xin_M_ffmem_mem_9__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3569 (
	.O(n2176),
	.A1(n2988),
	.A2(n2998),
	.B1B(n2988),
	.B2B(Mfifo_xin_M_ffmem_mem_9__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3570 (
	.O(n2177),
	.A1(n2988),
	.A2(n2997),
	.B1B(n2988),
	.B2B(Mfifo_xin_M_ffmem_mem_9__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3571 (
	.O(n2186),
	.A1(n2990),
	.A2(n3002),
	.B1B(n2990),
	.B2B(Mfifo_xin_M_ffmem_mem_11__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3572 (
	.O(n2187),
	.A1(n2990),
	.A2(n3001),
	.B1B(n2990),
	.B2B(Mfifo_xin_M_ffmem_mem_11__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3573 (
	.O(n2188),
	.A1(n2990),
	.A2(n3003),
	.B1B(n2990),
	.B2B(Mfifo_xin_M_ffmem_mem_11__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3574 (
	.O(n2189),
	.A1(n2990),
	.A2(n3005),
	.B1B(n2990),
	.B2B(Mfifo_xin_M_ffmem_mem_11__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3575 (
	.O(n2190),
	.A1(n2990),
	.A2(n3004),
	.B1B(n2990),
	.B2B(Mfifo_xin_M_ffmem_mem_11__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3576 (
	.O(n2191),
	.A1(n2990),
	.A2(n2999),
	.B1B(n2990),
	.B2B(Mfifo_xin_M_ffmem_mem_11__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3577 (
	.O(n2192),
	.A1(n2990),
	.A2(n2998),
	.B1B(n2990),
	.B2B(Mfifo_xin_M_ffmem_mem_11__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3578 (
	.O(n2206),
	.A1(n2991),
	.A2(n3004),
	.B1B(n2991),
	.B2B(Mfifo_xin_M_ffmem_mem_13__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3579 (
	.O(n2193),
	.A1(n2990),
	.A2(n2997),
	.B1B(n2990),
	.B2B(Mfifo_xin_M_ffmem_mem_11__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3580 (
	.O(n2208),
	.A1(n2991),
	.A2(n2998),
	.B1B(n2991),
	.B2B(Mfifo_xin_M_ffmem_mem_13__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3581 (
	.O(n2202),
	.A1(n2991),
	.A2(n3002),
	.B1B(n2991),
	.B2B(Mfifo_xin_M_ffmem_mem_13__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3582 (
	.O(n2203),
	.A1(n2991),
	.A2(n3001),
	.B1B(n2991),
	.B2B(Mfifo_xin_M_ffmem_mem_13__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3583 (
	.O(n2204),
	.A1(n2991),
	.A2(n3003),
	.B1B(n2991),
	.B2B(Mfifo_xin_M_ffmem_mem_13__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3584 (
	.O(n2205),
	.A1(n2991),
	.A2(n3005),
	.B1B(n2991),
	.B2B(Mfifo_xin_M_ffmem_mem_13__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3585 (
	.O(n2209),
	.A1(n2991),
	.A2(n2997),
	.B1B(n2991),
	.B2B(Mfifo_xin_M_ffmem_mem_13__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3586 (
	.O(n2207),
	.A1(n2991),
	.A2(n2999),
	.B1B(n2991),
	.B2B(Mfifo_xin_M_ffmem_mem_13__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3587 (
	.O(n2123),
	.A1(n2996),
	.A2(n3001),
	.B1B(n2996),
	.B2B(Mfifo_xin_M_ffmem_mem_3__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3588 (
	.O(n2112),
	.A1(n3006),
	.A2(n2998),
	.B1B(n3006),
	.B2B(Mfifo_xin_M_ffmem_mem_1__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3589 (
	.O(n2139),
	.A1(n3000),
	.A2(n3001),
	.B1B(n3000),
	.B2B(Mfifo_xin_M_ffmem_mem_5__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3590 (
	.O(n2138),
	.A1(n3000),
	.A2(n3002),
	.B1B(n3000),
	.B2B(Mfifo_xin_M_ffmem_mem_5__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3591 (
	.O(n2129),
	.A1(n2996),
	.A2(n2997),
	.B1B(n2996),
	.B2B(Mfifo_xin_M_ffmem_mem_3__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3592 (
	.O(n2128),
	.A1(n2996),
	.A2(n2998),
	.B1B(n2996),
	.B2B(Mfifo_xin_M_ffmem_mem_3__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3593 (
	.O(n2127),
	.A1(n2996),
	.A2(n2999),
	.B1B(n2996),
	.B2B(Mfifo_xin_M_ffmem_mem_3__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3594 (
	.O(n2126),
	.A1(n2996),
	.A2(n3004),
	.B1B(n2996),
	.B2B(Mfifo_xin_M_ffmem_mem_3__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3595 (
	.O(n2125),
	.A1(n2996),
	.A2(n3005),
	.B1B(n2996),
	.B2B(Mfifo_xin_M_ffmem_mem_3__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3596 (
	.O(n2124),
	.A1(n2996),
	.A2(n3003),
	.B1B(n2996),
	.B2B(Mfifo_xin_M_ffmem_mem_3__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3597 (
	.O(n2141),
	.A1(n3000),
	.A2(n3005),
	.B1B(n3000),
	.B2B(Mfifo_xin_M_ffmem_mem_5__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3598 (
	.O(n2122),
	.A1(n2996),
	.A2(n3002),
	.B1B(n2996),
	.B2B(Mfifo_xin_M_ffmem_mem_3__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3599 (
	.O(n2113),
	.A1(n3006),
	.A2(n2997),
	.B1B(n3006),
	.B2B(Mfifo_xin_M_ffmem_mem_1__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3600 (
	.O(n2145),
	.A1(n3000),
	.A2(n2997),
	.B1B(n3000),
	.B2B(Mfifo_xin_M_ffmem_mem_5__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3601 (
	.O(n2144),
	.A1(n3000),
	.A2(n2998),
	.B1B(n3000),
	.B2B(Mfifo_xin_M_ffmem_mem_5__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3602 (
	.O(n2143),
	.A1(n3000),
	.A2(n2999),
	.B1B(n3000),
	.B2B(Mfifo_xin_M_ffmem_mem_5__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3603 (
	.O(n2142),
	.A1(n3000),
	.A2(n3004),
	.B1B(n3000),
	.B2B(Mfifo_xin_M_ffmem_mem_5__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3604 (
	.O(n2111),
	.A1(n3006),
	.A2(n2999),
	.B1B(n3006),
	.B2B(Mfifo_xin_M_ffmem_mem_1__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3605 (
	.O(n2140),
	.A1(n3000),
	.A2(n3003),
	.B1B(n3000),
	.B2B(Mfifo_xin_M_ffmem_mem_5__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3606 (
	.O(n2107),
	.A1(n3006),
	.A2(n3001),
	.B1B(n3006),
	.B2B(Mfifo_xin_M_ffmem_mem_1__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3607 (
	.O(n2106),
	.A1(n3006),
	.A2(n3002),
	.B1B(n3006),
	.B2B(Mfifo_xin_M_ffmem_mem_1__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3608 (
	.O(n2108),
	.A1(n3006),
	.A2(n3003),
	.B1B(n3006),
	.B2B(Mfifo_xin_M_ffmem_mem_1__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3609 (
	.O(n2110),
	.A1(n3006),
	.A2(n3004),
	.B1B(n3006),
	.B2B(Mfifo_xin_M_ffmem_mem_1__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3610 (
	.O(n2109),
	.A1(n3006),
	.A2(n3005),
	.B1B(n3006),
	.B2B(Mfifo_xin_M_ffmem_mem_1__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3611 (
	.O(n2349),
	.A1(n3007),
	.A2(n3026),
	.B1B(n3007),
	.B2B(Mfifo_coe_M_ffmem_mem_14__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3612 (
	.O(n2347),
	.A1(n3007),
	.A2(n3021),
	.B1B(n3007),
	.B2B(Mfifo_coe_M_ffmem_mem_14__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3613 (
	.O(n2350),
	.A1(n3007),
	.A2(n3025),
	.B1B(n3007),
	.B2B(Mfifo_coe_M_ffmem_mem_14__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3614 (
	.O(n2346),
	.A1(n3007),
	.A2(n3023),
	.B1B(n3007),
	.B2B(Mfifo_coe_M_ffmem_mem_14__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3615 (
	.O(n2353),
	.A1(n3007),
	.A2(n3017),
	.B1B(n3007),
	.B2B(Mfifo_coe_M_ffmem_mem_14__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3616 (
	.O(n2351),
	.A1(n3007),
	.A2(n3027),
	.B1B(n3007),
	.B2B(Mfifo_coe_M_ffmem_mem_14__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3617 (
	.O(n2352),
	.A1(n3007),
	.A2(n3020),
	.B1B(n3007),
	.B2B(Mfifo_coe_M_ffmem_mem_14__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3618 (
	.O(n2348),
	.A1(n3007),
	.A2(n3019),
	.B1B(n3007),
	.B2B(Mfifo_coe_M_ffmem_mem_14__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U3619 (
	.O(n3009),
	.I1(n3008),
	.I2(n3016), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3620 (
	.O(n2321),
	.A1(n3009),
	.A2(n3017),
	.B1B(n3009),
	.B2B(Mfifo_coe_M_ffmem_mem_10__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3621 (
	.O(n2316),
	.A1(n3009),
	.A2(n3019),
	.B1B(n3009),
	.B2B(Mfifo_coe_M_ffmem_mem_10__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3622 (
	.O(n2317),
	.A1(n3009),
	.A2(n3026),
	.B1B(n3009),
	.B2B(Mfifo_coe_M_ffmem_mem_10__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U3623 (
	.O(n3010),
	.I1(n3008),
	.I2(n3013), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3624 (
	.O(n2298),
	.A1(n3010),
	.A2(n3023),
	.B1B(n3010),
	.B2B(Mfifo_coe_M_ffmem_mem_8__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U3625 (
	.O(n3011),
	.I1(n3008),
	.I2(n3014), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3626 (
	.O(n2332),
	.A1(n3011),
	.A2(n3019),
	.B1B(n3011),
	.B2B(Mfifo_coe_M_ffmem_mem_12__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3627 (
	.O(n2334),
	.A1(n3011),
	.A2(n3025),
	.B1B(n3011),
	.B2B(Mfifo_coe_M_ffmem_mem_12__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3628 (
	.O(n2303),
	.A1(n3010),
	.A2(n3027),
	.B1B(n3010),
	.B2B(Mfifo_coe_M_ffmem_mem_8__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3629 (
	.O(n2315),
	.A1(n3009),
	.A2(n3021),
	.B1B(n3009),
	.B2B(Mfifo_coe_M_ffmem_mem_10__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3630 (
	.O(n2305),
	.A1(n3010),
	.A2(n3017),
	.B1B(n3010),
	.B2B(Mfifo_coe_M_ffmem_mem_8__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3631 (
	.O(n2314),
	.A1(n3009),
	.A2(n3023),
	.B1B(n3009),
	.B2B(Mfifo_coe_M_ffmem_mem_10__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3632 (
	.O(n2330),
	.A1(n3011),
	.A2(n3023),
	.B1B(n3011),
	.B2B(Mfifo_coe_M_ffmem_mem_12__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3633 (
	.O(n2331),
	.A1(n3011),
	.A2(n3021),
	.B1B(n3011),
	.B2B(Mfifo_coe_M_ffmem_mem_12__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3634 (
	.O(n2299),
	.A1(n3010),
	.A2(n3021),
	.B1B(n3010),
	.B2B(Mfifo_coe_M_ffmem_mem_8__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3635 (
	.O(n2318),
	.A1(n3009),
	.A2(n3025),
	.B1B(n3009),
	.B2B(Mfifo_coe_M_ffmem_mem_10__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3636 (
	.O(n2319),
	.A1(n3009),
	.A2(n3027),
	.B1B(n3009),
	.B2B(Mfifo_coe_M_ffmem_mem_10__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3637 (
	.O(n2320),
	.A1(n3009),
	.A2(n3020),
	.B1B(n3009),
	.B2B(Mfifo_coe_M_ffmem_mem_10__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3638 (
	.O(n2336),
	.A1(n3011),
	.A2(n3020),
	.B1B(n3011),
	.B2B(Mfifo_coe_M_ffmem_mem_12__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3639 (
	.O(n2304),
	.A1(n3010),
	.A2(n3020),
	.B1B(n3010),
	.B2B(Mfifo_coe_M_ffmem_mem_8__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3640 (
	.O(n2335),
	.A1(n3011),
	.A2(n3027),
	.B1B(n3011),
	.B2B(Mfifo_coe_M_ffmem_mem_12__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3641 (
	.O(n2302),
	.A1(n3010),
	.A2(n3025),
	.B1B(n3010),
	.B2B(Mfifo_coe_M_ffmem_mem_8__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3642 (
	.O(n2300),
	.A1(n3010),
	.A2(n3019),
	.B1B(n3010),
	.B2B(Mfifo_coe_M_ffmem_mem_8__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3643 (
	.O(n2301),
	.A1(n3010),
	.A2(n3026),
	.B1B(n3010),
	.B2B(Mfifo_coe_M_ffmem_mem_8__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3644 (
	.O(n2333),
	.A1(n3011),
	.A2(n3026),
	.B1B(n3011),
	.B2B(Mfifo_coe_M_ffmem_mem_12__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3645 (
	.O(n2337),
	.A1(n3011),
	.A2(n3017),
	.B1B(n3011),
	.B2B(Mfifo_coe_M_ffmem_mem_12__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3646 (
	.O(n2241),
	.A1(n3022),
	.A2(n3017),
	.B1B(n3022),
	.B2B(Mfifo_coe_M_ffmem_mem_0__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3647 (
	.O(n2237),
	.A1(n3022),
	.A2(n3026),
	.B1B(n3022),
	.B2B(Mfifo_coe_M_ffmem_mem_0__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3648 (
	.O(n2238),
	.A1(n3022),
	.A2(n3025),
	.B1B(n3022),
	.B2B(Mfifo_coe_M_ffmem_mem_0__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3649 (
	.O(n2239),
	.A1(n3022),
	.A2(n3027),
	.B1B(n3022),
	.B2B(Mfifo_coe_M_ffmem_mem_0__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3650 (
	.O(n2283),
	.A1(n3024),
	.A2(n3021),
	.B1B(n3024),
	.B2B(Mfifo_coe_M_ffmem_mem_6__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3651 (
	.O(n2284),
	.A1(n3024),
	.A2(n3019),
	.B1B(n3024),
	.B2B(Mfifo_coe_M_ffmem_mem_6__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3652 (
	.O(n2240),
	.A1(n3022),
	.A2(n3020),
	.B1B(n3022),
	.B2B(Mfifo_coe_M_ffmem_mem_0__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3653 (
	.O(n2289),
	.A1(n3024),
	.A2(n3017),
	.B1B(n3024),
	.B2B(Mfifo_coe_M_ffmem_mem_6__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3654 (
	.O(n2288),
	.A1(n3024),
	.A2(n3020),
	.B1B(n3024),
	.B2B(Mfifo_coe_M_ffmem_mem_6__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3655 (
	.O(n2287),
	.A1(n3024),
	.A2(n3027),
	.B1B(n3024),
	.B2B(Mfifo_coe_M_ffmem_mem_6__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3656 (
	.O(n2286),
	.A1(n3024),
	.A2(n3025),
	.B1B(n3024),
	.B2B(Mfifo_coe_M_ffmem_mem_6__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3657 (
	.O(n2267),
	.A1(n3028),
	.A2(n3021),
	.B1B(n3028),
	.B2B(Mfifo_coe_M_ffmem_mem_4__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3658 (
	.O(n2268),
	.A1(n3028),
	.A2(n3019),
	.B1B(n3028),
	.B2B(Mfifo_coe_M_ffmem_mem_4__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3659 (
	.O(n2250),
	.A1(n3018),
	.A2(n3023),
	.B1B(n3018),
	.B2B(Mfifo_coe_M_ffmem_mem_2__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3660 (
	.O(n2234),
	.A1(n3022),
	.A2(n3023),
	.B1B(n3022),
	.B2B(Mfifo_coe_M_ffmem_mem_0__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3661 (
	.O(n2251),
	.A1(n3018),
	.A2(n3021),
	.B1B(n3018),
	.B2B(Mfifo_coe_M_ffmem_mem_2__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3662 (
	.O(n2252),
	.A1(n3018),
	.A2(n3019),
	.B1B(n3018),
	.B2B(Mfifo_coe_M_ffmem_mem_2__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3663 (
	.O(n2253),
	.A1(n3018),
	.A2(n3026),
	.B1B(n3018),
	.B2B(Mfifo_coe_M_ffmem_mem_2__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3664 (
	.O(n2254),
	.A1(n3018),
	.A2(n3025),
	.B1B(n3018),
	.B2B(Mfifo_coe_M_ffmem_mem_2__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3665 (
	.O(n2255),
	.A1(n3018),
	.A2(n3027),
	.B1B(n3018),
	.B2B(Mfifo_coe_M_ffmem_mem_2__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3666 (
	.O(n2256),
	.A1(n3018),
	.A2(n3020),
	.B1B(n3018),
	.B2B(Mfifo_coe_M_ffmem_mem_2__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3667 (
	.O(n2273),
	.A1(n3028),
	.A2(n3017),
	.B1B(n3028),
	.B2B(Mfifo_coe_M_ffmem_mem_4__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3668 (
	.O(n2257),
	.A1(n3018),
	.A2(n3017),
	.B1B(n3018),
	.B2B(Mfifo_coe_M_ffmem_mem_2__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3669 (
	.O(n2266),
	.A1(n3028),
	.A2(n3023),
	.B1B(n3028),
	.B2B(Mfifo_coe_M_ffmem_mem_4__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3670 (
	.O(n2236),
	.A1(n3022),
	.A2(n3019),
	.B1B(n3022),
	.B2B(Mfifo_coe_M_ffmem_mem_0__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3671 (
	.O(n2272),
	.A1(n3028),
	.A2(n3020),
	.B1B(n3028),
	.B2B(Mfifo_coe_M_ffmem_mem_4__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3672 (
	.O(n2235),
	.A1(n3022),
	.A2(n3021),
	.B1B(n3022),
	.B2B(Mfifo_coe_M_ffmem_mem_0__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3673 (
	.O(n2282),
	.A1(n3024),
	.A2(n3023),
	.B1B(n3024),
	.B2B(Mfifo_coe_M_ffmem_mem_6__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3674 (
	.O(n2285),
	.A1(n3024),
	.A2(n3026),
	.B1B(n3024),
	.B2B(Mfifo_coe_M_ffmem_mem_6__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3675 (
	.O(n2270),
	.A1(n3028),
	.A2(n3025),
	.B1B(n3028),
	.B2B(Mfifo_coe_M_ffmem_mem_4__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3676 (
	.O(n2269),
	.A1(n3028),
	.A2(n3026),
	.B1B(n3028),
	.B2B(Mfifo_coe_M_ffmem_mem_4__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3677 (
	.O(n2271),
	.A1(n3028),
	.A2(n3027),
	.B1B(n3028),
	.B2B(Mfifo_coe_M_ffmem_mem_4__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3678 (
	.O(Mfifo_psum_M_rptr_rbinnext[0]),
	.A1(n3032),
	.B1(n3030),
	.B2(n3029), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3679 (
	.O(Mfifo_psum_M_rptr_rbinnext[1]),
	.A1(n3037),
	.B1(Mfifo_psum_raddr[1]),
	.B2(n3032), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3680 (
	.O(Mfifo_psum_M_rptr_rgraynext[0]),
	.A1(Mfifo_psum_M_rptr_rbinnext[0]),
	.A2(Mfifo_psum_raddr[1]),
	.B1B(Mfifo_psum_M_rptr_rbinnext[0]),
	.B2B(Mfifo_psum_M_rptr_rbinnext[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U3681 (
	.O(n3217),
	.B2(n3031),
	.I1(n3032), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3682 (
	.O(Mfifo_psum_M_rptr_rbinnext[4]),
	.A1(Mfifo_psum_rptr[4]),
	.A2(n3217),
	.B1B(Mfifo_psum_rptr[4]),
	.B2B(n3217), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3683 (
	.O(n3218),
	.I1(Mfifo_psum_raddr[3]),
	.I2(n3033), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3684 (
	.O(n3034),
	.I1(Mfifo_psum_M_rptr_rbinnext[4]),
	.I2(n3218), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3685 (
	.O(Mfifo_psum_M_rptr_rgraynext[3]),
	.A1(n3034),
	.B1(n3218),
	.B2(Mfifo_psum_rptr[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3686 (
	.O(Mfifo_psum_M_rptr_rgraynext[2]),
	.A1(Mfifo_psum_raddr[3]),
	.A2(n3035),
	.B1B(Mfifo_psum_raddr[3]),
	.B2B(n3035), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3687 (
	.O(Mfifo_psum_M_rptr_rgraynext[1]),
	.A1(n3037),
	.A2(n3036),
	.B1B(n3036),
	.B2B(n3037), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3688 (
	.O(n3047),
	.I(Mfifo_psum_M_rptr_rgraynext[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3689 (
	.O(n3040),
	.I(Mfifo_psum_M_rptr_rgraynext[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3690 (
	.O(n3039),
	.I(Mfifo_psum_M_rptr_rgraynext[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3691 (
	.O(n3038),
	.A1(n3040),
	.A2(Mfifo_psum_rq2_wptr[3]),
	.B1(n3039),
	.B2(Mfifo_psum_rq2_wptr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3692 (
	.O(n3045),
	.A1(n3038),
	.B1(n3040),
	.B2(Mfifo_psum_rq2_wptr[3]),
	.C1(Mfifo_psum_rq2_wptr[2]),
	.C2(n3039), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3693 (
	.O(n3043),
	.I(Mfifo_psum_M_rptr_rbinnext[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3694 (
	.O(n3042),
	.I(Mfifo_psum_M_rptr_rgraynext[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3695 (
	.O(n3041),
	.A1(n3043),
	.A2(Mfifo_psum_rq2_wptr[4]),
	.B1(Mfifo_psum_rq2_wptr[1]),
	.B2(n3042), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3696 (
	.O(n3044),
	.A1(n3041),
	.B1(n3043),
	.B2(Mfifo_psum_rq2_wptr[4]),
	.C1(n3042),
	.C2(Mfifo_psum_rq2_wptr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3697 (
	.O(n3046),
	.A1(n3045),
	.B1(n3044),
	.C1(n3047),
	.C2(Mfifo_psum_rq2_wptr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3698 (
	.O(Mfifo_psum_M_rptr_rempty_val),
	.A1(n3046),
	.B1(n3047),
	.B2(Mfifo_psum_rq2_wptr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3699 (
	.O(n3211),
	.I1(n3049),
	.I2(n3048), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI21B1X05AR9 U3700 (
	.O(Mfifo_xin_M_wptr_wbinnext[3]),
	.A1(n3211),
	.A2(n3052),
	.B1B(n3050), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3701 (
	.O(Mfifo_xin_M_wptr_wbinnext[4]),
	.A1(Mfifo_xin_wptr[4]),
	.A2(n3051),
	.B1B(n3051),
	.B2B(Mfifo_xin_wptr[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3702 (
	.O(Mfifo_xin_M_wptr_wgraynext[3]),
	.A1(Mfifo_xin_M_wptr_wbinnext[3]),
	.A2(Mfifo_xin_wptr[4]),
	.B1B(Mfifo_xin_M_wptr_wbinnext[3]),
	.B2B(Mfifo_xin_M_wptr_wbinnext[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3703 (
	.O(n3210),
	.A1(Mfifo_xin_waddr[2]),
	.B1(Mfifo_xin_waddr[1]),
	.B2(n3213), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3704 (
	.O(Mfifo_xin_M_wptr_wgraynext[2]),
	.A1(n3210),
	.A2(n3052),
	.B1B(n3210),
	.B2B(n3052), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3705 (
	.O(Mfifo_xin_M_wptr_wgraynext[1]),
	.A1(Mfifo_xin_waddr[2]),
	.A2(n3053),
	.B1B(Mfifo_xin_waddr[2]),
	.B2B(n3053), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3706 (
	.O(n3212),
	.I1(Mfifo_xin_waddr[0]),
	.I2(n3054), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3707 (
	.O(Mfifo_xin_M_wptr_wgraynext[0]),
	.A1(n3212),
	.A2(n3055),
	.B1B(n3212),
	.B2B(n3055), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3708 (
	.O(n3057),
	.I(Mfifo_xin_M_wptr_wgraynext[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3709 (
	.O(n3056),
	.A1(Mfifo_xin_M_wptr_wbinnext[4]),
	.A2(Mfifo_xin_wq2_rptr[4]),
	.B1(Mfifo_xin_wq2_rptr[2]),
	.B2(n3057), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3710 (
	.O(n3062),
	.A1(n3056),
	.B1(Mfifo_xin_M_wptr_wbinnext[4]),
	.B2(Mfifo_xin_wq2_rptr[4]),
	.C1(n3057),
	.C2(Mfifo_xin_wq2_rptr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3711 (
	.O(n3060),
	.I(Mfifo_xin_M_wptr_wgraynext[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3712 (
	.O(n3059),
	.I(Mfifo_xin_M_wptr_wgraynext[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3713 (
	.O(n3058),
	.A1(n3060),
	.A2(Mfifo_xin_wq2_rptr[1]),
	.B1(n3059),
	.B2(Mfifo_xin_wq2_rptr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3714 (
	.O(n3061),
	.A1(n3058),
	.B1(n3060),
	.B2(Mfifo_xin_wq2_rptr[1]),
	.C1(Mfifo_xin_wq2_rptr[0]),
	.C2(n3059), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3715 (
	.O(n3063),
	.A1(n3062),
	.B1(n3061),
	.C1(Mfifo_xin_wq2_rptr[3]),
	.C2(Mfifo_xin_M_wptr_wgraynext[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3716 (
	.O(Mfifo_xin_M_wptr_wfull_val),
	.A1(n3063),
	.B1(Mfifo_xin_wq2_rptr[3]),
	.B2(Mfifo_xin_M_wptr_wgraynext[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3717 (
	.O(Mfifo_coe_M_wptr_wbinnext[4]),
	.A1(n3064),
	.A2(Mfifo_coe_wptr[4]),
	.B1B(Mfifo_coe_wptr[4]),
	.B2B(n3064), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3718 (
	.O(n3220),
	.A1(Mfifo_coe_waddr[2]),
	.B1(Mfifo_coe_waddr[1]),
	.B2(n3222), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3719 (
	.O(Mfifo_coe_M_wptr_wgraynext[2]),
	.A1(n3220),
	.A2(n3068),
	.B1B(n3220),
	.B2B(n3068), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3720 (
	.O(n3219),
	.I1(n3066),
	.I2(n3065), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI21B1X05AR9 U3721 (
	.O(Mfifo_coe_M_wptr_wbinnext[3]),
	.A1(n3219),
	.A2(n3068),
	.B1B(n3067), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3722 (
	.O(Mfifo_coe_M_wptr_wgraynext[3]),
	.A1(Mfifo_coe_M_wptr_wbinnext[3]),
	.A2(Mfifo_coe_wptr[4]),
	.B1B(Mfifo_coe_M_wptr_wbinnext[3]),
	.B2B(Mfifo_coe_M_wptr_wbinnext[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3723 (
	.O(Mfifo_coe_M_wptr_wgraynext[1]),
	.A1(Mfifo_coe_waddr[2]),
	.A2(n3069),
	.B1B(Mfifo_coe_waddr[2]),
	.B2B(n3069), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3724 (
	.O(n3221),
	.I1(Mfifo_coe_waddr[0]),
	.I2(n3070), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3725 (
	.O(Mfifo_coe_M_wptr_wgraynext[0]),
	.A1(n3221),
	.A2(n3071),
	.B1B(n3221),
	.B2B(n3071), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3726 (
	.O(n3073),
	.I(Mfifo_coe_M_wptr_wgraynext[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3727 (
	.O(n3072),
	.A1(n3073),
	.A2(Mfifo_coe_wq2_rptr[2]),
	.B1(Mfifo_coe_wq2_rptr[3]),
	.B2(Mfifo_coe_M_wptr_wgraynext[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3728 (
	.O(n3078),
	.A1(n3072),
	.B1(n3073),
	.B2(Mfifo_coe_wq2_rptr[2]),
	.C1(Mfifo_coe_M_wptr_wgraynext[3]),
	.C2(Mfifo_coe_wq2_rptr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3729 (
	.O(n3076),
	.I(Mfifo_coe_M_wptr_wgraynext[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3730 (
	.O(n3075),
	.I(Mfifo_coe_M_wptr_wgraynext[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3731 (
	.O(n3074),
	.A1(n3076),
	.A2(Mfifo_coe_wq2_rptr[1]),
	.B1(n3075),
	.B2(Mfifo_coe_wq2_rptr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3732 (
	.O(n3077),
	.A1(n3074),
	.B1(n3076),
	.B2(Mfifo_coe_wq2_rptr[1]),
	.C1(Mfifo_coe_wq2_rptr[0]),
	.C2(n3075), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3733 (
	.O(n3079),
	.A1(n3078),
	.B1(n3077),
	.C1(Mfifo_coe_M_wptr_wbinnext[4]),
	.C2(Mfifo_coe_wq2_rptr[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3734 (
	.O(Mfifo_coe_M_wptr_wfull_val),
	.A1(n3079),
	.B1(Mfifo_coe_M_wptr_wbinnext[4]),
	.B2(Mfifo_coe_wq2_rptr[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3735 (
	.O(n1386),
	.A1(n3829),
	.A2(n3113),
	.B1B(n3829),
	.B2B(int_H[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3736 (
	.O(n1389),
	.A1(n3829),
	.A2(n3514),
	.B1B(n3829),
	.B2B(int_W[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3737 (
	.O(n1390),
	.A1(n3829),
	.A2(n3523),
	.B1B(n3829),
	.B2B(int_W[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3738 (
	.O(n3251),
	.I(Mcntl_flag), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3739 (
	.O(n3320),
	.I(n3317), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3740 (
	.O(n2376),
	.A1(n3320),
	.B1(n3080),
	.B2(n3251), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3741 (
	.O(n3081),
	.I1(n3827),
	.I2(int_ky[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3742 (
	.O(n1391),
	.A1(n3081),
	.B1(n3827),
	.B2(n3082), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3743 (
	.O(n3288),
	.I(Mcntl_Mcntldata_kx_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3744 (
	.O(n3083),
	.I1(n3827),
	.I2(int_kx[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3745 (
	.O(n1382),
	.A1(n3083),
	.B1(n3827),
	.B2(n3288), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3746 (
	.O(n3086),
	.I1(count_k[0]),
	.I2(count_k[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3747 (
	.O(n3084),
	.A1(count_k[0]),
	.A2(count_k[1]),
	.B1(count_k[2]),
	.B2(n3086), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3748 (
	.O(n2389),
	.I1(n3084),
	.I2(n3839), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3749 (
	.O(n3085),
	.I(count_k[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3750 (
	.O(n2387),
	.A1(n3839),
	.B1(n3086),
	.B2(n3085), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2X05AR9 U3751 (
	.O(n3174),
	.I1(int_ky[0]),
	.I2(n3827), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI21B1X05AR9 U3752 (
	.O(n1392),
	.A1(n3827),
	.A2(n3087),
	.B1B(n3174), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3753 (
	.O(n3098),
	.I1(Mcntl_Mcntldata_c_W_d4[1]),
	.I2(n3109), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3754 (
	.O(n3094),
	.A1(n3106),
	.B1(n3091),
	.B2(n3512), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3755 (
	.O(n3088),
	.A1(Mcntl_Mcntldata_c_W_d4[0]),
	.A2(n3098),
	.B1(n3094),
	.B2(n3310), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI13X05AR9 U3756 (
	.O(n3089),
	.A1(n3088),
	.B1(n3091),
	.B2(n3090),
	.B3(n3310), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3757 (
	.O(n3524),
	.I(Mcntl_Mcntldata_c_W_d4[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3758 (
	.O(n3107),
	.I(n3096), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3759 (
	.O(n2083),
	.A1(n3096),
	.A2(n3089),
	.B1(n3524),
	.B2(n3107), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3760 (
	.O(n3092),
	.I1(n3091),
	.I2(n3090), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3761 (
	.O(n3095),
	.A1(n3094),
	.A2(n3093),
	.B1(n3312),
	.B2(n3092), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3762 (
	.O(n3097),
	.A1(n3096),
	.A2(n3095),
	.B1(Mcntl_Mcntldata_c_W_d4[1]),
	.B2(n3107), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3763 (
	.O(n2089),
	.A1(n3097),
	.B1(n3524),
	.B2(n3098), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3764 (
	.O(n3239),
	.I1(psum_wfull),
	.I2(n3099), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3765 (
	.O(n3242),
	.I(n3239), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI13X05AR9 U3766 (
	.O(n3102),
	.A1(Mcntl_Mcntl_current_state[2]),
	.B1(n3101),
	.B2(n3100),
	.B3(n3242), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3767 (
	.O(n2394),
	.I1(n3102),
	.I2(n3320), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U3768 (
	.O(n3105),
	.I1(Mcntl_Mcntldata_c_cin[0]),
	.I2(c_cout[3]),
	.I3(n3274), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U3769 (
	.O(n3103),
	.I1(c_cout[0]),
	.I2(c_cout[1]),
	.I3(c_cout[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR3B2X05AR9 U3770 (
	.O(n3231),
	.B2(n3105),
	.B3(n3103),
	.I1(Mcntl_Mcntldata_c_cin[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR4X05AR9 U3771 (
	.O(n3268),
	.I1(c_cout[0]),
	.I2(c_cout[1]),
	.I3(c_cout[2]),
	.I4(n3267), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3772 (
	.O(n3275),
	.I1(n3105),
	.I2(n3268), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12B2X05AR9 U3773 (
	.O(n2378),
	.A1(n3829),
	.B1B(Mcntl_Mcntldata_c_cin[1]),
	.B2B(n3275), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12B2X05AR9 U3774 (
	.O(n3519),
	.A1(n3106),
	.B1B(n3108),
	.B2B(n3107), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3775 (
	.O(n3518),
	.A1(n3519),
	.B1(Mcntl_Mcntldata_c_x_cin[0]),
	.B2(n3109), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3776 (
	.O(n2082),
	.A1(n3110),
	.B1(n3518),
	.B2(n3111), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3777 (
	.O(n3115),
	.I(Mcntl_Mcntldata_c_x_H[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI21B1X05AR9 U3778 (
	.O(n3184),
	.A1(Mcntl_Mcntldata_x_H_reg[0]),
	.A2(Mcntl_Mcntldata_ky_reg[0]),
	.B1B(n3112), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI222X05AR9 U3779 (
	.O(n3114),
	.A1(n3121),
	.A2(n3113),
	.B1(n3115),
	.B2(n3122),
	.C1(n3184),
	.C2(n3125), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3780 (
	.O(n2084),
	.A1(n3129),
	.A2(n3115),
	.B1(n3114),
	.B2(n3126), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3781 (
	.O(n3299),
	.A1(n3116),
	.B1(n3120),
	.B2(n3117), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3782 (
	.O(n3124),
	.I(n3299), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3783 (
	.O(n3123),
	.A1(n3118),
	.B1(n3119),
	.B2(n3128), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI222X05AR9 U3784 (
	.O(n3127),
	.A1(n3125),
	.A2(n3124),
	.B1(n3123),
	.B2(n3122),
	.C1(n3121),
	.C2(n3120), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3785 (
	.O(n2086),
	.A1(n3129),
	.A2(n3128),
	.B1(n3127),
	.B2(n3126), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3786 (
	.O(Mfifo_xin_M_rptr_rgraynext[3]),
	.A1(Mfifo_xin_rptr[4]),
	.A2(n3130),
	.B1B(Mfifo_xin_rptr[4]),
	.B2B(n3130), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3787 (
	.O(Mfifo_xin_M_rptr_rbinnext[4]),
	.A1(Mfifo_xin_rptr[4]),
	.A2(n3131),
	.B1B(Mfifo_xin_rptr[4]),
	.B2B(n3131), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3788 (
	.O(Mfifo_xin_M_rptr_rgraynext[2]),
	.A1(n3132),
	.A2(n3419),
	.B1B(n3132),
	.B2B(n3419), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3789 (
	.O(Mfifo_xin_M_rptr_rgraynext[1]),
	.A1(Mfifo_xin_raddr[2]),
	.A2(n3133),
	.B1B(Mfifo_xin_raddr[2]),
	.B2B(n3133), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3790 (
	.O(n3216),
	.I1(Mfifo_xin_M_rptr_N1),
	.I2(Mfifo_xin_raddr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3791 (
	.O(Mfifo_xin_M_rptr_rgraynext[0]),
	.A1(n3216),
	.A2(n3418),
	.B1B(n3216),
	.B2B(n3418), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3792 (
	.O(n3143),
	.I(Mfifo_xin_M_rptr_rgraynext[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3793 (
	.O(n3136),
	.I(Mfifo_xin_M_rptr_rbinnext[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3794 (
	.O(n3135),
	.I(Mfifo_xin_M_rptr_rgraynext[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3795 (
	.O(n3134),
	.A1(n3136),
	.A2(Mfifo_xin_rq2_wptr[4]),
	.B1(n3135),
	.B2(Mfifo_xin_rq2_wptr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3796 (
	.O(n3141),
	.A1(n3134),
	.B1(n3136),
	.B2(Mfifo_xin_rq2_wptr[4]),
	.C1(Mfifo_xin_rq2_wptr[2]),
	.C2(n3135), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3797 (
	.O(n3139),
	.I(Mfifo_xin_M_rptr_rgraynext[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3798 (
	.O(n3138),
	.I(Mfifo_xin_M_rptr_rgraynext[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3799 (
	.O(n3137),
	.A1(n3139),
	.A2(Mfifo_xin_rq2_wptr[1]),
	.B1(n3138),
	.B2(Mfifo_xin_rq2_wptr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3800 (
	.O(n3140),
	.A1(n3137),
	.B1(n3139),
	.B2(Mfifo_xin_rq2_wptr[1]),
	.C1(Mfifo_xin_rq2_wptr[0]),
	.C2(n3138), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3801 (
	.O(n3142),
	.A1(n3141),
	.B1(n3140),
	.C1(n3143),
	.C2(Mfifo_xin_rq2_wptr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3802 (
	.O(Mfifo_xin_M_rptr_rempty_val),
	.A1(n3142),
	.B1(n3143),
	.B2(Mfifo_xin_rq2_wptr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2B1X05AR9 U3803 (
	.O(n3273),
	.B2(n3268),
	.I1(c_cout[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3804 (
	.O(n3271),
	.I1(n3829),
	.I2(n3273), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3805 (
	.O(n3249),
	.I1(xen4),
	.I2(n3271), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3806 (
	.O(n3166),
	.I1(n3173),
	.I2(n3267), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3807 (
	.O(n3167),
	.I1(c_kx[1]),
	.I2(n3166), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3808 (
	.O(n3168),
	.I(n3166), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3809 (
	.O(n3245),
	.A1(n3164),
	.B1(n3168),
	.B2(n3144), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3810 (
	.O(n3145),
	.A1(n3827),
	.A2(int_kx[0]),
	.B1(Mcntl_Mcntldata_kx_reg[0]),
	.B2(n3245), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3811 (
	.O(n3146),
	.A1(n3145),
	.B1(c_kx[0]),
	.B2(n3167), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3812 (
	.O(n2379),
	.A1(n3249),
	.A2(n3224),
	.B1B(n3249),
	.B2B(n3146), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3813 (
	.O(n3279),
	.I(n3277), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3814 (
	.O(n3149),
	.I1(Mcntl_Mcntldata_c_p_cout[1]),
	.I2(n3279), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3815 (
	.O(n3148),
	.I(Mcntl_Mcntldata_c_p_cout[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3816 (
	.O(n3291),
	.I1(n3280),
	.I2(n3147), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3817 (
	.O(n3189),
	.I(n3291), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3818 (
	.O(n2373),
	.A1(n3189),
	.B1(n3149),
	.B2(n3148), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3819 (
	.O(Mfifo_coe_M_rptr_rbinnext[4]),
	.A1(Mfifo_coe_rptr[4]),
	.A2(n3150),
	.B1B(Mfifo_coe_rptr[4]),
	.B2B(n3150), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3820 (
	.O(Mfifo_coe_M_rptr_rgraynext[2]),
	.A1(Mfifo_coe_raddr[3]),
	.A2(n3151),
	.B1B(Mfifo_coe_raddr[3]),
	.B2B(n3151), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3821 (
	.O(Mfifo_coe_M_rptr_rgraynext[3]),
	.A1(Mfifo_coe_rptr[4]),
	.A2(n3152),
	.B1B(Mfifo_coe_rptr[4]),
	.B2B(n3152), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3822 (
	.O(Mfifo_coe_M_rptr_rgraynext[1]),
	.A1(n3153),
	.A2(n3325),
	.B1B(n3153),
	.B2B(n3325), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3823 (
	.O(n3223),
	.I1(Mfifo_coe_M_rptr_N1),
	.I2(Mfifo_coe_raddr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3824 (
	.O(Mfifo_coe_M_rptr_rgraynext[0]),
	.A1(n3223),
	.A2(n3326),
	.B1B(n3223),
	.B2B(n3326), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3825 (
	.O(n3163),
	.I(Mfifo_coe_M_rptr_rbinnext[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3826 (
	.O(n3156),
	.I(Mfifo_coe_M_rptr_rgraynext[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3827 (
	.O(n3155),
	.I(Mfifo_coe_M_rptr_rgraynext[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3828 (
	.O(n3154),
	.A1(n3156),
	.A2(Mfifo_coe_rq2_wptr[2]),
	.B1(n3155),
	.B2(Mfifo_coe_rq2_wptr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3829 (
	.O(n3161),
	.A1(n3154),
	.B1(n3156),
	.B2(Mfifo_coe_rq2_wptr[2]),
	.C1(Mfifo_coe_rq2_wptr[3]),
	.C2(n3155), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3830 (
	.O(n3159),
	.I(Mfifo_coe_M_rptr_rgraynext[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3831 (
	.O(n3158),
	.I(Mfifo_coe_M_rptr_rgraynext[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3832 (
	.O(n3157),
	.A1(n3159),
	.A2(Mfifo_coe_rq2_wptr[1]),
	.B1(n3158),
	.B2(Mfifo_coe_rq2_wptr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3833 (
	.O(n3160),
	.A1(n3157),
	.B1(n3159),
	.B2(Mfifo_coe_rq2_wptr[1]),
	.C1(Mfifo_coe_rq2_wptr[0]),
	.C2(n3158), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3834 (
	.O(n3162),
	.A1(n3161),
	.B1(n3160),
	.C1(n3163),
	.C2(Mfifo_coe_rq2_wptr[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3835 (
	.O(Mfifo_coe_M_rptr_rempty_val),
	.A1(n3162),
	.B1(n3163),
	.B2(Mfifo_coe_rq2_wptr[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3836 (
	.O(n3176),
	.A1(n3164),
	.B1(n3165),
	.B2(n3267), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3837 (
	.O(n3171),
	.A1(n3827),
	.A2(int_ky[1]),
	.B1(Mcntl_Mcntldata_ky_reg[1]),
	.B2(n3176), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3838 (
	.O(n3247),
	.A1(n3249),
	.B1(c_kx[0]),
	.B2(n3166), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3839 (
	.O(n3177),
	.I1(n3247),
	.I2(n3167), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3840 (
	.O(n3169),
	.I1(n3168),
	.I2(n3178), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3841 (
	.O(n3170),
	.A1(c_ky[1]),
	.B1(n3169),
	.B2(n3177), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3842 (
	.O(n2386),
	.A1(n3170),
	.B1(n3171),
	.B2(n3177), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3843 (
	.O(n3180),
	.I(n3177), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U3844 (
	.O(n3175),
	.A1(n3172),
	.B1(c_ky[0]),
	.C1(n3173),
	.C2(n3267), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U3845 (
	.O(n3179),
	.A1(n3175),
	.B1(n3174),
	.C1(Mcntl_Mcntldata_ky_reg[0]),
	.C2(n3176), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3846 (
	.O(n2385),
	.A1(n3180),
	.A2(n3179),
	.B1(n3178),
	.B2(n3177), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3847 (
	.O(n3284),
	.A1(n3291),
	.B1(n3263),
	.B2(n3190), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U3848 (
	.O(n3182),
	.I1(n3320),
	.I2(n3839),
	.I3(n3284), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3849 (
	.O(n3302),
	.A1(n3188),
	.B1(n3181),
	.B2(n3311), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3850 (
	.O(n3301),
	.I1(n3182),
	.I2(n3302), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3851 (
	.O(n3229),
	.I1(Mcntl_Mcntldata_c_p_wd4[1]),
	.I2(Mcntl_Mcntldata_c_p_wd4[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3852 (
	.O(n3304),
	.A1(n3182),
	.B1(n3229),
	.B2(n3839), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3853 (
	.O(n3306),
	.I1(n3183),
	.I2(n3320), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3854 (
	.O(n3185),
	.A1(Mcntl_Mcntldata_c_p_H[0]),
	.A2(n3304),
	.B1(n3184),
	.B2(n3306), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3855 (
	.O(n2369),
	.A1(n3185),
	.B1(Mcntl_Mcntldata_c_p_H[0]),
	.B2(n3301), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3856 (
	.O(n3286),
	.I1(Mcntl_Mcntldata_x_W_reg[0]),
	.I2(n3288), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3857 (
	.O(n3257),
	.I1(n3187),
	.I2(n3186), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA12X05AR9 U3858 (
	.O(n3192),
	.A1(n3257),
	.B1(n3187),
	.B2(n3186), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR4X05AR9 U3859 (
	.O(n3281),
	.I1(sel_reg[0]),
	.I2(n3190),
	.I3(n3189),
	.I4(n3188), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3860 (
	.O(n3537),
	.I(sel_reg[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3861 (
	.O(n3282),
	.I1(n3281),
	.I2(n3537), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3862 (
	.O(n3262),
	.I1(Mcntl_Mcntldata_c_p_W[2]),
	.I2(n3282), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI13X05AR9 U3863 (
	.O(n3191),
	.A1(n3262),
	.B1(Mcntl_Mcntldata_c_p_W[2]),
	.B2(n3280),
	.B3(n3282), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3864 (
	.O(n2371),
	.A1(n3191),
	.B1(n3192),
	.B2(n3284), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3865 (
	.O(n3550),
	.I(n3193), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3866 (
	.O(n3214),
	.A1(Mfifo_psum_waddr[2]),
	.B1(n3550),
	.B2(Mfifo_psum_waddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3867 (
	.O(n3543),
	.I(Mfifo_psum_waddr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3868 (
	.O(Mfifo_psum_M_wptr_wgraynext[2]),
	.A1(n3214),
	.A2(n3543),
	.B1B(n3214),
	.B2B(n3543), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3869 (
	.O(n3535),
	.I1(Mfifo_psum_waddr[2]),
	.I2(Mfifo_psum_waddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3870 (
	.O(Mfifo_psum_M_wptr_wgraynext[1]),
	.A1(Mfifo_psum_waddr[2]),
	.A2(n3194),
	.B1(n3535),
	.B2(n3193), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3871 (
	.O(n3215),
	.I1(n3549),
	.I2(Mfifo_psum_waddr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3872 (
	.O(Mfifo_psum_M_wptr_wgraynext[0]),
	.A1(n3215),
	.A2(n3544),
	.B1B(n3215),
	.B2B(n3544), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3873 (
	.O(n3196),
	.I(Mfifo_psum_M_wptr_wgraynext[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3874 (
	.O(n3195),
	.A1(Mfifo_psum_M_wptr_wbinnext[4]),
	.A2(Mfifo_psum_wq2_rptr[4]),
	.B1(n3196),
	.B2(Mfifo_psum_wq2_rptr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3875 (
	.O(n3201),
	.A1(n3195),
	.B1(Mfifo_psum_M_wptr_wbinnext[4]),
	.B2(Mfifo_psum_wq2_rptr[4]),
	.C1(Mfifo_psum_wq2_rptr[2]),
	.C2(n3196), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3876 (
	.O(n3199),
	.I(Mfifo_psum_M_wptr_wgraynext[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3877 (
	.O(n3198),
	.I(Mfifo_psum_M_wptr_wgraynext[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3878 (
	.O(n3197),
	.A1(n3199),
	.A2(Mfifo_psum_wq2_rptr[1]),
	.B1(n3198),
	.B2(Mfifo_psum_wq2_rptr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI122X05AR9 U3879 (
	.O(n3200),
	.A1(n3197),
	.B1(n3199),
	.B2(Mfifo_psum_wq2_rptr[1]),
	.C1(Mfifo_psum_wq2_rptr[0]),
	.C2(n3198), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3880 (
	.O(n3202),
	.A1(n3201),
	.B1(n3200),
	.C1(Mfifo_psum_wq2_rptr[3]),
	.C2(Mfifo_psum_M_wptr_wgraynext[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3881 (
	.O(Mfifo_psum_M_wptr_wfull_val),
	.A1(n3202),
	.B1(Mfifo_psum_wq2_rptr[3]),
	.B2(Mfifo_psum_M_wptr_wgraynext[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3882 (
	.O(n3203),
	.A1(n3288),
	.B1(c_kx[0]),
	.B2(n3246), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U3883 (
	.O(n2396),
	.A1(n3203),
	.B1(n3246),
	.B2(Mcntl_Mcntldata_kx_reg[1]),
	.C1(c_kx[0]),
	.C2(n3288), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3884 (
	.O(DP_OP_1207J5_130_8771_n12),
	.I(Mcntl_Mcntldata_N453), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   XOR2X05AR9 U3885 (
	.O(n3204),
	.I1(x_addr[6]),
	.I2(C2_Z_0), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3886 (
	.O(n3206),
	.I(n3205), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO22X05AR9 U3887 (
	.O(n3832),
	.A1(n3207),
	.A2(n2916),
	.B1(x_addr[6]),
	.B2(n3206), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3889 (
	.O(Mfifo_xin_M_wptr_wbinnext[2]),
	.I1(n3211),
	.I2(n3210), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3890 (
	.O(Mfifo_xin_M_wptr_wbinnext[0]),
	.I1(n3213),
	.I2(n3212), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3891 (
	.O(Mfifo_psum_M_wptr_wbinnext[2]),
	.I1(n3547),
	.I2(n3214), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3892 (
	.O(Mfifo_psum_M_wptr_wbinnext[0]),
	.I1(n3550),
	.I2(n3215), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3893 (
	.O(Mfifo_xin_M_rptr_rbinnext[0]),
	.I1(n3510),
	.I2(n3216), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3894 (
	.O(Mfifo_psum_M_rptr_rbinnext[3]),
	.I1(n3218),
	.I2(n3217), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3895 (
	.O(Mfifo_coe_M_wptr_wbinnext[2]),
	.I1(n3220),
	.I2(n3219), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3896 (
	.O(Mfifo_coe_M_wptr_wbinnext[0]),
	.I1(n3222),
	.I2(n3221), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3897 (
	.O(Mfifo_coe_M_rptr_rbinnext[0]),
	.I1(n3416),
	.I2(n3223), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3898 (
	.O(n3227),
	.I(n2396), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3899 (
	.O(n3226),
	.A1(n3246),
	.B1(c_kx[0]),
	.B2(n3288), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U3900 (
	.O(n3225),
	.A1(c_kx[1]),
	.B1(n3224),
	.C1(Mcntl_Mcntldata_kx_reg[1]),
	.C2(Mcntl_Mcntldata_kx_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3901 (
	.O(n2397),
	.A1(Mcntl_Mcntldata_kx_reg[1]),
	.A2(n3227),
	.B1(n3226),
	.B2(n3225), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3902 (
	.O(n3230),
	.I(n3529), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3903 (
	.O(n3528),
	.I1(n3229),
	.I2(n3228), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3904 (
	.O(n3237),
	.A1(int_end_read),
	.B1(n3230),
	.B2(n3528), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI13X05AR9 U3905 (
	.O(n3234),
	.A1(n3252),
	.B1(n3233),
	.B2(n3232),
	.B3(n3231), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U3906 (
	.O(n3236),
	.A1(n3263),
	.B1(n3827),
	.C1(n3235),
	.C2(n3234), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3907 (
	.O(n2395),
	.A1(n3237),
	.B1(n3236),
	.C1(n3239),
	.C2(n3238), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3908 (
	.O(n3526),
	.I(n3240), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3909 (
	.O(n3243),
	.I1(Mcntl_Mcntl_current_state[2]),
	.I2(Mcntl_Mcntl_current_state[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3910 (
	.O(n3244),
	.A1(Mcntl_Mcntl_current_state[1]),
	.B1(n3241),
	.C1(n3243),
	.C2(n3242), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3911 (
	.O(n2393),
	.A1(n3526),
	.B1(n3244),
	.C1(n3529),
	.C2(n3528), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3912 (
	.O(n3248),
	.A1(n3827),
	.A2(int_kx[1]),
	.B1(Mcntl_Mcntldata_kx_reg[1]),
	.B2(n3245), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U3913 (
	.O(n2392),
	.A1(n3249),
	.A2(n3248),
	.B1(n3247),
	.B2(n3246), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3914 (
	.O(n3253),
	.A1(n3250),
	.B1(Mcntl_Mcntldata_count[1]),
	.C1(Mcntl_Mcntl_current_state[0]),
	.C2(n3251), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3915 (
	.O(n3256),
	.I(Mcntl_Mcntldata_count[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2B1X05AR9 U3916 (
	.O(n3254),
	.B2(n3251),
	.I1(n3252), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U3917 (
	.O(n2391),
	.A1(n3254),
	.B1(Mcntl_Mcntldata_count[0]),
	.B2(n3253),
	.C1(n3256),
	.C2(n3255), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U3918 (
	.O(n2390),
	.A1(n3254),
	.B1(n3530),
	.B2(n3256),
	.C1(n3530),
	.C2(n3255), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3919 (
	.O(n3261),
	.I(Mcntl_Mcntldata_c_p_W[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3920 (
	.O(n3259),
	.I(n3257), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3921 (
	.O(n3287),
	.I(n3284), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U3922 (
	.O(n3260),
	.A1(n3287),
	.B1(Mcntl_Mcntldata_x_W_reg[3]),
	.B2(n3259),
	.C1(n3258),
	.C2(n3257), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI13X05AR9 U3923 (
	.O(n2384),
	.A1(n3260),
	.B1(n3263),
	.B2(n3262),
	.B3(n3261), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3924 (
	.O(n3264),
	.I1(n3267),
	.I2(c_cout[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO112X05AR9 U3925 (
	.O(n2383),
	.A1(n3827),
	.B1(n3264),
	.C1(n3267),
	.C2(c_cout[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3926 (
	.O(n3266),
	.I(n3264), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3927 (
	.O(n3265),
	.I(c_cout[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U3928 (
	.O(n2382),
	.A1(n3829),
	.B1(c_cout[1]),
	.B2(n3266),
	.C1(n3265),
	.C2(n3264), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X05AR9 U3929 (
	.O(n3270),
	.I1(c_cout[0]),
	.I2(c_cout[1]),
	.I3(n3267), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3930 (
	.O(n3269),
	.I(c_cout[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3931 (
	.O(n3272),
	.I(n3268), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3932 (
	.O(n2381),
	.A1(n3272),
	.B1(n3829),
	.C1(n3270),
	.C2(n3269), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO12X05AR9 U3933 (
	.O(n2380),
	.A1(n3271),
	.B1(c_cout[3]),
	.B2(n3272), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3934 (
	.O(n3276),
	.A1(Mcntl_Mcntldata_c_cin[0]),
	.B1(n3274),
	.B2(n3273), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U3935 (
	.O(n2377),
	.I1(n3829),
	.I2(n3276),
	.I3(n3275), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3936 (
	.O(n3278),
	.I(Mcntl_Mcntldata_c_p_cout[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U3937 (
	.O(n2375),
	.A1(n3280),
	.B1(Mcntl_Mcntldata_c_p_cout[1]),
	.B2(n3279),
	.C1(n3278),
	.C2(n3277), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3938 (
	.O(n2374),
	.A1(n3280),
	.B1(n3279),
	.C1(n3549),
	.C2(n3805), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3939 (
	.O(n3290),
	.I(n3281), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3940 (
	.O(n3285),
	.I1(sel_reg[1]),
	.I2(n3290), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U3941 (
	.O(n2372),
	.A1(n3282),
	.B1(n3287),
	.B2(n3285),
	.C1(n3284),
	.C2(n3283), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3942 (
	.O(n3536),
	.I(sel_reg[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3943 (
	.O(n3289),
	.A1(n3287),
	.B1(n3286),
	.C1(Mcntl_Mcntldata_x_W_reg[0]),
	.C2(n3288), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3944 (
	.O(n2370),
	.A1(n3290),
	.B1(n3289),
	.C1(n3291),
	.C2(n3536), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3945 (
	.O(n3296),
	.I(n3292), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3946 (
	.O(n3300),
	.I(n3306), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3947 (
	.O(n3294),
	.I(Mcntl_Mcntldata_c_p_H[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3948 (
	.O(n3293),
	.A1(n3304),
	.B1(Mcntl_Mcntldata_c_p_H[0]),
	.B2(n3302), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI222X05AR9 U3949 (
	.O(n2368),
	.A1(n3301),
	.A2(n3296),
	.B1(n3300),
	.B2(n3295),
	.C1(n3294),
	.C2(n3293), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U3950 (
	.O(n3297),
	.A1(n3304),
	.B1(n3296),
	.B2(n3302), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI222X05AR9 U3951 (
	.O(n2367),
	.A1(n3301),
	.A2(n3303),
	.B1(n3300),
	.B2(n3299),
	.C1(n3298),
	.C2(n3297), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U3952 (
	.O(n3305),
	.A1(Mcntl_Mcntldata_c_p_H[3]),
	.B1(n3304),
	.B2(n3303),
	.C1(n3304),
	.C2(n3302), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12B2X05AR9 U3953 (
	.O(n2366),
	.A1(n3305),
	.B1B(n3307),
	.B2B(n3306), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U3954 (
	.O(n3309),
	.I1(Mcntl_Mcntldata_c_p_wd4[0]),
	.I2(n3320),
	.I3(n3839), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U3955 (
	.O(n3308),
	.A1(n3316),
	.B1(Mcntl_Mcntldata_c_p_wd4[1]),
	.B2(n3310), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3956 (
	.O(n2365),
	.A1(n3309),
	.B1(n3308),
	.C1(n3310),
	.C2(n3320), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U3957 (
	.O(n3314),
	.A1(n3317),
	.A2(n3313),
	.B1B(n3312),
	.B2B(n3311), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI13X05AR9 U3958 (
	.O(n2364),
	.A1(n3314),
	.B1(n3317),
	.B2(n3316),
	.B3(n3315), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3959 (
	.O(n3318),
	.I(Mcntl_Mcntldata_c_p_cin[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U3960 (
	.O(n3323),
	.I1(n3319),
	.I2(n3318), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U3961 (
	.O(n2363),
	.A1(n3320),
	.B1(n3323),
	.C1(n3319),
	.C2(n3318), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3962 (
	.O(n3322),
	.I(Mcntl_Mcntldata_c_p_cin[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U3963 (
	.O(n3321),
	.I(n3323), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U3964 (
	.O(n2362),
	.A1(n3320),
	.B1(Mcntl_Mcntldata_c_p_cin[1]),
	.B2(n3323),
	.C1(n3322),
	.C2(n3321), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U3965 (
	.O(n3404),
	.I1(Mfifo_coe_raddr[1]),
	.I2(Mfifo_coe_raddr[3]),
	.I3(n3325), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U3966 (
	.O(n3402),
	.I1(Mfifo_coe_raddr[1]),
	.I2(n3324),
	.I3(n3325), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3967 (
	.O(n3330),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_5__1_),
	.B1(n3402),
	.B2(Mfifo_coe_M_ffmem_mem_13__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U3968 (
	.O(n3401),
	.I1(Mfifo_coe_raddr[1]),
	.I2(Mfifo_coe_raddr[2]),
	.I3(n3324), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U3969 (
	.O(n3408),
	.I1(Mfifo_coe_raddr[2]),
	.I2(n3324),
	.I3(n3326), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3970 (
	.O(n3329),
	.A1(n3401),
	.A2(Mfifo_coe_M_ffmem_mem_9__1_),
	.B1(n3408),
	.B2(Mfifo_coe_M_ffmem_mem_11__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U3971 (
	.O(n3403),
	.I1(Mfifo_coe_raddr[3]),
	.I2(n3326),
	.I3(n3325), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U3972 (
	.O(n3407),
	.I1(Mfifo_coe_raddr[1]),
	.I2(Mfifo_coe_raddr[3]),
	.I3(Mfifo_coe_raddr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3973 (
	.O(n3328),
	.A1(n3403),
	.A2(Mfifo_coe_M_ffmem_mem_7__1_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_1__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U3974 (
	.O(n3405),
	.I1(Mfifo_coe_raddr[3]),
	.I2(Mfifo_coe_raddr[2]),
	.I3(n3326), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3975 (
	.O(n3327),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_15__1_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_3__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3976 (
	.O(n3336),
	.I1(n3330),
	.I2(n3329),
	.I3(n3328),
	.I4(n3327), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3977 (
	.O(n3334),
	.A1(n3403),
	.A2(Mfifo_coe_M_ffmem_mem_6__1_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_2__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3978 (
	.O(n3333),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_4__1_),
	.B1(n3402),
	.B2(Mfifo_coe_M_ffmem_mem_12__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3979 (
	.O(n3332),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_14__1_),
	.B1(n3408),
	.B2(Mfifo_coe_M_ffmem_mem_10__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3980 (
	.O(n3331),
	.A1(n3401),
	.A2(Mfifo_coe_M_ffmem_mem_8__1_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_0__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3981 (
	.O(n3335),
	.I1(n3334),
	.I2(n3333),
	.I3(n3332),
	.I4(n3331), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U3982 (
	.O(n3413),
	.I1(Mfifo_coe_raddr[0]),
	.I2(n3415), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U3983 (
	.O(n2233),
	.A1(n3336),
	.A2(n3416),
	.B1(n3415),
	.B2(int_coe[1]),
	.C1(n3335),
	.C2(n3413), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3984 (
	.O(n3340),
	.A1(n3401),
	.A2(Mfifo_coe_M_ffmem_mem_9__2_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_3__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3985 (
	.O(n3339),
	.A1(n3402),
	.A2(Mfifo_coe_M_ffmem_mem_13__2_),
	.B1(n3403),
	.B2(Mfifo_coe_M_ffmem_mem_7__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3986 (
	.O(n3338),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_15__2_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_1__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3987 (
	.O(n3337),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_5__2_),
	.B1(n3408),
	.B2(Mfifo_coe_M_ffmem_mem_11__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3988 (
	.O(n3346),
	.I1(n3340),
	.I2(n3339),
	.I3(n3338),
	.I4(n3337), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3989 (
	.O(n3344),
	.A1(n3402),
	.A2(Mfifo_coe_M_ffmem_mem_12__2_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_0__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3990 (
	.O(n3343),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_14__2_),
	.B1(n3408),
	.B2(Mfifo_coe_M_ffmem_mem_10__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3991 (
	.O(n3342),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_4__2_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_2__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3992 (
	.O(n3341),
	.A1(n3401),
	.A2(Mfifo_coe_M_ffmem_mem_8__2_),
	.B1(n3403),
	.B2(Mfifo_coe_M_ffmem_mem_6__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3993 (
	.O(n3345),
	.I1(n3344),
	.I2(n3343),
	.I3(n3342),
	.I4(n3341), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U3994 (
	.O(n2232),
	.A1(n3346),
	.A2(n3416),
	.B1(n3415),
	.B2(int_coe[2]),
	.C1(n3345),
	.C2(n3413), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3995 (
	.O(n3350),
	.A1(n3408),
	.A2(Mfifo_coe_M_ffmem_mem_11__3_),
	.B1(n3403),
	.B2(Mfifo_coe_M_ffmem_mem_7__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3996 (
	.O(n3349),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_15__3_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_3__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3997 (
	.O(n3348),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_5__3_),
	.B1(n3401),
	.B2(Mfifo_coe_M_ffmem_mem_9__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U3998 (
	.O(n3347),
	.A1(n3402),
	.A2(Mfifo_coe_M_ffmem_mem_13__3_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_1__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U3999 (
	.O(n3356),
	.I1(n3350),
	.I2(n3349),
	.I3(n3348),
	.I4(n3347), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4000 (
	.O(n3354),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_14__3_),
	.B1(n3408),
	.B2(Mfifo_coe_M_ffmem_mem_10__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4001 (
	.O(n3353),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_4__3_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_0__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4002 (
	.O(n3352),
	.A1(n3402),
	.A2(Mfifo_coe_M_ffmem_mem_12__3_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_2__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4003 (
	.O(n3351),
	.A1(n3401),
	.A2(Mfifo_coe_M_ffmem_mem_8__3_),
	.B1(n3403),
	.B2(Mfifo_coe_M_ffmem_mem_6__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4004 (
	.O(n3355),
	.I1(n3354),
	.I2(n3353),
	.I3(n3352),
	.I4(n3351), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4005 (
	.O(n2231),
	.A1(n3356),
	.A2(n3416),
	.B1(n3415),
	.B2(int_coe[3]),
	.C1(n3355),
	.C2(n3413), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4006 (
	.O(n3360),
	.A1(n3402),
	.A2(Mfifo_coe_M_ffmem_mem_13__4_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_3__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4007 (
	.O(n3359),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_15__4_),
	.B1(n3403),
	.B2(Mfifo_coe_M_ffmem_mem_7__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4008 (
	.O(n3358),
	.A1(n3408),
	.A2(Mfifo_coe_M_ffmem_mem_11__4_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_1__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4009 (
	.O(n3357),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_5__4_),
	.B1(n3401),
	.B2(Mfifo_coe_M_ffmem_mem_9__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4010 (
	.O(n3366),
	.I1(n3360),
	.I2(n3359),
	.I3(n3358),
	.I4(n3357), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4011 (
	.O(n3364),
	.A1(n3403),
	.A2(Mfifo_coe_M_ffmem_mem_6__4_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_0__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4012 (
	.O(n3363),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_14__4_),
	.B1(n3408),
	.B2(Mfifo_coe_M_ffmem_mem_10__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4013 (
	.O(n3362),
	.A1(n3402),
	.A2(Mfifo_coe_M_ffmem_mem_12__4_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_2__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4014 (
	.O(n3361),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_4__4_),
	.B1(n3401),
	.B2(Mfifo_coe_M_ffmem_mem_8__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4015 (
	.O(n3365),
	.I1(n3364),
	.I2(n3363),
	.I3(n3362),
	.I4(n3361), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4016 (
	.O(n2230),
	.A1(n3366),
	.A2(n3416),
	.B1(n3415),
	.B2(int_coe[4]),
	.C1(n3365),
	.C2(n3413), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4017 (
	.O(n3370),
	.A1(n3401),
	.A2(Mfifo_coe_M_ffmem_mem_9__5_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_3__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4018 (
	.O(n3369),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_5__5_),
	.B1(n3408),
	.B2(Mfifo_coe_M_ffmem_mem_11__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4019 (
	.O(n3368),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_15__5_),
	.B1(n3402),
	.B2(Mfifo_coe_M_ffmem_mem_13__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4020 (
	.O(n3367),
	.A1(n3403),
	.A2(Mfifo_coe_M_ffmem_mem_7__5_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_1__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4021 (
	.O(n3376),
	.I1(n3370),
	.I2(n3369),
	.I3(n3368),
	.I4(n3367), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4022 (
	.O(n3374),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_4__5_),
	.B1(n3401),
	.B2(Mfifo_coe_M_ffmem_mem_8__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4023 (
	.O(n3373),
	.A1(n3403),
	.A2(Mfifo_coe_M_ffmem_mem_6__5_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_0__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4024 (
	.O(n3372),
	.A1(n3408),
	.A2(Mfifo_coe_M_ffmem_mem_10__5_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_2__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4025 (
	.O(n3371),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_14__5_),
	.B1(n3402),
	.B2(Mfifo_coe_M_ffmem_mem_12__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4026 (
	.O(n3375),
	.I1(n3374),
	.I2(n3373),
	.I3(n3372),
	.I4(n3371), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4027 (
	.O(n2229),
	.A1(n3376),
	.A2(n3416),
	.B1(n3415),
	.B2(int_coe[5]),
	.C1(n3375),
	.C2(n3413), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4028 (
	.O(n3380),
	.A1(n3408),
	.A2(Mfifo_coe_M_ffmem_mem_11__6_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_1__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4029 (
	.O(n3379),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_5__6_),
	.B1(n3403),
	.B2(Mfifo_coe_M_ffmem_mem_7__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4030 (
	.O(n3378),
	.A1(n3402),
	.A2(Mfifo_coe_M_ffmem_mem_13__6_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_3__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4031 (
	.O(n3377),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_15__6_),
	.B1(n3401),
	.B2(Mfifo_coe_M_ffmem_mem_9__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4032 (
	.O(n3386),
	.I1(n3380),
	.I2(n3379),
	.I3(n3378),
	.I4(n3377), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4033 (
	.O(n3384),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_14__6_),
	.B1(n3403),
	.B2(Mfifo_coe_M_ffmem_mem_6__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4034 (
	.O(n3383),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_4__6_),
	.B1(n3402),
	.B2(Mfifo_coe_M_ffmem_mem_12__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4035 (
	.O(n3382),
	.A1(n3408),
	.A2(Mfifo_coe_M_ffmem_mem_10__6_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_2__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4036 (
	.O(n3381),
	.A1(n3401),
	.A2(Mfifo_coe_M_ffmem_mem_8__6_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_0__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4037 (
	.O(n3385),
	.I1(n3384),
	.I2(n3383),
	.I3(n3382),
	.I4(n3381), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4038 (
	.O(n2228),
	.A1(n3386),
	.A2(n3416),
	.B1(n3415),
	.B2(int_coe[6]),
	.C1(n3385),
	.C2(n3413), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4039 (
	.O(n3390),
	.A1(n3402),
	.A2(Mfifo_coe_M_ffmem_mem_13__7_),
	.B1(n3408),
	.B2(Mfifo_coe_M_ffmem_mem_11__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4040 (
	.O(n3389),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_15__7_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_3__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4041 (
	.O(n3388),
	.A1(n3401),
	.A2(Mfifo_coe_M_ffmem_mem_9__7_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_1__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4042 (
	.O(n3387),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_5__7_),
	.B1(n3403),
	.B2(Mfifo_coe_M_ffmem_mem_7__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4043 (
	.O(n3396),
	.I1(n3390),
	.I2(n3389),
	.I3(n3388),
	.I4(n3387), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4044 (
	.O(n3394),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_4__7_),
	.B1(n3408),
	.B2(Mfifo_coe_M_ffmem_mem_10__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4045 (
	.O(n3393),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_14__7_),
	.B1(n3403),
	.B2(Mfifo_coe_M_ffmem_mem_6__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4046 (
	.O(n3392),
	.A1(n3402),
	.A2(Mfifo_coe_M_ffmem_mem_12__7_),
	.B1(n3401),
	.B2(Mfifo_coe_M_ffmem_mem_8__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4047 (
	.O(n3391),
	.A1(n3407),
	.A2(Mfifo_coe_M_ffmem_mem_0__7_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_2__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4048 (
	.O(n3395),
	.I1(n3394),
	.I2(n3393),
	.I3(n3392),
	.I4(n3391), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4049 (
	.O(n2227),
	.A1(n3396),
	.A2(n3416),
	.B1(n3415),
	.B2(int_coe[7]),
	.C1(n3395),
	.C2(n3413), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4050 (
	.O(n3400),
	.A1(n3407),
	.A2(Mfifo_coe_M_ffmem_mem_1__0_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_3__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4051 (
	.O(n3399),
	.A1(n3402),
	.A2(Mfifo_coe_M_ffmem_mem_13__0_),
	.B1(n3403),
	.B2(Mfifo_coe_M_ffmem_mem_7__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4052 (
	.O(n3398),
	.A1(n3401),
	.A2(Mfifo_coe_M_ffmem_mem_9__0_),
	.B1(n3408),
	.B2(Mfifo_coe_M_ffmem_mem_11__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4053 (
	.O(n3397),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_15__0_),
	.B1(n3404),
	.B2(Mfifo_coe_M_ffmem_mem_5__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4054 (
	.O(n3417),
	.I1(n3400),
	.I2(n3399),
	.I3(n3398),
	.I4(n3397), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4055 (
	.O(n3412),
	.A1(n3402),
	.A2(Mfifo_coe_M_ffmem_mem_12__0_),
	.B1(n3401),
	.B2(Mfifo_coe_M_ffmem_mem_8__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4056 (
	.O(n3411),
	.A1(n3404),
	.A2(Mfifo_coe_M_ffmem_mem_4__0_),
	.B1(n3403),
	.B2(Mfifo_coe_M_ffmem_mem_6__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4057 (
	.O(n3410),
	.A1(n3406),
	.A2(Mfifo_coe_M_ffmem_mem_14__0_),
	.B1(n3405),
	.B2(Mfifo_coe_M_ffmem_mem_2__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4058 (
	.O(n3409),
	.A1(n3408),
	.A2(Mfifo_coe_M_ffmem_mem_10__0_),
	.B1(n3407),
	.B2(Mfifo_coe_M_ffmem_mem_0__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4059 (
	.O(n3414),
	.I1(n3412),
	.I2(n3411),
	.I3(n3410),
	.I4(n3409), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4060 (
	.O(n2226),
	.A1(n3417),
	.A2(n3416),
	.B1(n3415),
	.B2(int_coe[0]),
	.C1(n3414),
	.C2(n3413), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U4061 (
	.O(n3496),
	.I1(Mfifo_xin_raddr[3]),
	.I2(Mfifo_xin_raddr[2]),
	.I3(Mfifo_xin_raddr[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U4062 (
	.O(n3502),
	.I1(Mfifo_xin_raddr[1]),
	.I2(n3420),
	.I3(n3419), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4063 (
	.O(n3424),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_1__1_),
	.B1(n3502),
	.B2(Mfifo_xin_M_ffmem_mem_13__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U4064 (
	.O(n3497),
	.I1(Mfifo_xin_raddr[3]),
	.I2(n3420),
	.I3(n3418), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U4065 (
	.O(n3495),
	.I1(Mfifo_xin_raddr[2]),
	.I2(n3419),
	.I3(n3418), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4066 (
	.O(n3423),
	.A1(n3497),
	.A2(Mfifo_xin_M_ffmem_mem_7__1_),
	.B1(n3495),
	.B2(Mfifo_xin_M_ffmem_mem_11__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U4067 (
	.O(n3500),
	.I1(Mfifo_xin_raddr[3]),
	.I2(Mfifo_xin_raddr[2]),
	.I3(n3418), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4068 (
	.O(n3422),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_15__1_),
	.B1(n3500),
	.B2(Mfifo_xin_M_ffmem_mem_3__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U4069 (
	.O(n3501),
	.I1(Mfifo_xin_raddr[2]),
	.I2(Mfifo_xin_raddr[1]),
	.I3(n3419), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U4070 (
	.O(n3499),
	.I1(Mfifo_xin_raddr[3]),
	.I2(Mfifo_xin_raddr[1]),
	.I3(n3420), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4071 (
	.O(n3421),
	.A1(n3501),
	.A2(Mfifo_xin_M_ffmem_mem_9__1_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_5__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4072 (
	.O(n3430),
	.I1(n3424),
	.I2(n3423),
	.I3(n3422),
	.I4(n3421), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4073 (
	.O(n3509),
	.I(Mfifo_xin_M_rptr_N1), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4074 (
	.O(n3428),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_0__1_),
	.B1(n3495),
	.B2(Mfifo_xin_M_ffmem_mem_10__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4075 (
	.O(n3427),
	.A1(n3502),
	.A2(Mfifo_xin_M_ffmem_mem_12__1_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_8__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4076 (
	.O(n3426),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_14__1_),
	.B1(n3500),
	.B2(Mfifo_xin_M_ffmem_mem_2__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4077 (
	.O(n3425),
	.A1(n3497),
	.A2(Mfifo_xin_M_ffmem_mem_6__1_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_4__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4078 (
	.O(n3429),
	.I1(n3428),
	.I2(n3427),
	.I3(n3426),
	.I4(n3425), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U4079 (
	.O(n3507),
	.I1(Mfifo_xin_raddr[0]),
	.I2(n3509), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4080 (
	.O(n2097),
	.A1(n3430),
	.A2(n3510),
	.B1(n3509),
	.B2(int_xin[1]),
	.C1(n3429),
	.C2(n3507), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4081 (
	.O(n3434),
	.A1(n3501),
	.A2(Mfifo_xin_M_ffmem_mem_9__2_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_5__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4082 (
	.O(n3433),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_15__2_),
	.B1(n3495),
	.B2(Mfifo_xin_M_ffmem_mem_11__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4083 (
	.O(n3432),
	.A1(n3497),
	.A2(Mfifo_xin_M_ffmem_mem_7__2_),
	.B1(n3500),
	.B2(Mfifo_xin_M_ffmem_mem_3__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4084 (
	.O(n3431),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_1__2_),
	.B1(n3502),
	.B2(Mfifo_xin_M_ffmem_mem_13__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4085 (
	.O(n3440),
	.I1(n3434),
	.I2(n3433),
	.I3(n3432),
	.I4(n3431), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4086 (
	.O(n3438),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_14__2_),
	.B1(n3500),
	.B2(Mfifo_xin_M_ffmem_mem_2__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4087 (
	.O(n3437),
	.A1(n3502),
	.A2(Mfifo_xin_M_ffmem_mem_12__2_),
	.B1(n3497),
	.B2(Mfifo_xin_M_ffmem_mem_6__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4088 (
	.O(n3436),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_0__2_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_4__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4089 (
	.O(n3435),
	.A1(n3495),
	.A2(Mfifo_xin_M_ffmem_mem_10__2_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_8__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4090 (
	.O(n3439),
	.I1(n3438),
	.I2(n3437),
	.I3(n3436),
	.I4(n3435), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4091 (
	.O(n2096),
	.A1(n3440),
	.A2(n3510),
	.B1(n3509),
	.B2(int_xin[2]),
	.C1(n3439),
	.C2(n3507), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4092 (
	.O(n3444),
	.A1(n3497),
	.A2(Mfifo_xin_M_ffmem_mem_7__3_),
	.B1(n3500),
	.B2(Mfifo_xin_M_ffmem_mem_3__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4093 (
	.O(n3443),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_15__3_),
	.B1(n3496),
	.B2(Mfifo_xin_M_ffmem_mem_1__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4094 (
	.O(n3442),
	.A1(n3502),
	.A2(Mfifo_xin_M_ffmem_mem_13__3_),
	.B1(n3495),
	.B2(Mfifo_xin_M_ffmem_mem_11__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4095 (
	.O(n3441),
	.A1(n3501),
	.A2(Mfifo_xin_M_ffmem_mem_9__3_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_5__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4096 (
	.O(n3450),
	.I1(n3444),
	.I2(n3443),
	.I3(n3442),
	.I4(n3441), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4097 (
	.O(n3448),
	.A1(n3500),
	.A2(Mfifo_xin_M_ffmem_mem_2__3_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_8__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4098 (
	.O(n3447),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_14__3_),
	.B1(n3502),
	.B2(Mfifo_xin_M_ffmem_mem_12__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4099 (
	.O(n3446),
	.A1(n3497),
	.A2(Mfifo_xin_M_ffmem_mem_6__3_),
	.B1(n3495),
	.B2(Mfifo_xin_M_ffmem_mem_10__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4100 (
	.O(n3445),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_0__3_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_4__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4101 (
	.O(n3449),
	.I1(n3448),
	.I2(n3447),
	.I3(n3446),
	.I4(n3445), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4102 (
	.O(n2095),
	.A1(n3450),
	.A2(n3510),
	.B1(n3509),
	.B2(int_xin[3]),
	.C1(n3449),
	.C2(n3507), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4103 (
	.O(n3454),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_1__4_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_9__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4104 (
	.O(n3453),
	.A1(n3500),
	.A2(Mfifo_xin_M_ffmem_mem_3__4_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_5__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4105 (
	.O(n3452),
	.A1(n3502),
	.A2(Mfifo_xin_M_ffmem_mem_13__4_),
	.B1(n3497),
	.B2(Mfifo_xin_M_ffmem_mem_7__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4106 (
	.O(n3451),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_15__4_),
	.B1(n3495),
	.B2(Mfifo_xin_M_ffmem_mem_11__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4107 (
	.O(n3460),
	.I1(n3454),
	.I2(n3453),
	.I3(n3452),
	.I4(n3451), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4108 (
	.O(n3458),
	.A1(n3502),
	.A2(Mfifo_xin_M_ffmem_mem_12__4_),
	.B1(n3500),
	.B2(Mfifo_xin_M_ffmem_mem_2__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4109 (
	.O(n3457),
	.A1(n3497),
	.A2(Mfifo_xin_M_ffmem_mem_6__4_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_4__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4110 (
	.O(n3456),
	.A1(n3495),
	.A2(Mfifo_xin_M_ffmem_mem_10__4_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_8__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4111 (
	.O(n3455),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_14__4_),
	.B1(n3496),
	.B2(Mfifo_xin_M_ffmem_mem_0__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4112 (
	.O(n3459),
	.I1(n3458),
	.I2(n3457),
	.I3(n3456),
	.I4(n3455), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4113 (
	.O(n2094),
	.A1(n3460),
	.A2(n3510),
	.B1(n3509),
	.B2(int_xin[4]),
	.C1(n3459),
	.C2(n3507), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4114 (
	.O(n3464),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_15__5_),
	.B1(n3495),
	.B2(Mfifo_xin_M_ffmem_mem_11__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4115 (
	.O(n3463),
	.A1(n3502),
	.A2(Mfifo_xin_M_ffmem_mem_13__5_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_5__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4116 (
	.O(n3462),
	.A1(n3497),
	.A2(Mfifo_xin_M_ffmem_mem_7__5_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_9__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4117 (
	.O(n3461),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_1__5_),
	.B1(n3500),
	.B2(Mfifo_xin_M_ffmem_mem_3__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4118 (
	.O(n3470),
	.I1(n3464),
	.I2(n3463),
	.I3(n3462),
	.I4(n3461), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4119 (
	.O(n3468),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_14__5_),
	.B1(n3497),
	.B2(Mfifo_xin_M_ffmem_mem_6__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4120 (
	.O(n3467),
	.A1(n3500),
	.A2(Mfifo_xin_M_ffmem_mem_2__5_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_4__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4121 (
	.O(n3466),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_0__5_),
	.B1(n3502),
	.B2(Mfifo_xin_M_ffmem_mem_12__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4122 (
	.O(n3465),
	.A1(n3495),
	.A2(Mfifo_xin_M_ffmem_mem_10__5_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_8__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4123 (
	.O(n3469),
	.I1(n3468),
	.I2(n3467),
	.I3(n3466),
	.I4(n3465), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4124 (
	.O(n2093),
	.A1(n3470),
	.A2(n3510),
	.B1(n3509),
	.B2(int_xin[5]),
	.C1(n3469),
	.C2(n3507), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4125 (
	.O(n3474),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_1__6_),
	.B1(n3495),
	.B2(Mfifo_xin_M_ffmem_mem_11__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4126 (
	.O(n3473),
	.A1(n3502),
	.A2(Mfifo_xin_M_ffmem_mem_13__6_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_9__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4127 (
	.O(n3472),
	.A1(n3497),
	.A2(Mfifo_xin_M_ffmem_mem_7__6_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_5__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4128 (
	.O(n3471),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_15__6_),
	.B1(n3500),
	.B2(Mfifo_xin_M_ffmem_mem_3__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4129 (
	.O(n3480),
	.I1(n3474),
	.I2(n3473),
	.I3(n3472),
	.I4(n3471), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4130 (
	.O(n3478),
	.A1(n3495),
	.A2(Mfifo_xin_M_ffmem_mem_10__6_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_4__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4131 (
	.O(n3477),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_14__6_),
	.B1(n3502),
	.B2(Mfifo_xin_M_ffmem_mem_12__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4132 (
	.O(n3476),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_0__6_),
	.B1(n3500),
	.B2(Mfifo_xin_M_ffmem_mem_2__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4133 (
	.O(n3475),
	.A1(n3497),
	.A2(Mfifo_xin_M_ffmem_mem_6__6_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_8__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4134 (
	.O(n3479),
	.I1(n3478),
	.I2(n3477),
	.I3(n3476),
	.I4(n3475), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4135 (
	.O(n2092),
	.A1(n3480),
	.A2(n3510),
	.B1(n3509),
	.B2(int_xin[6]),
	.C1(n3479),
	.C2(n3507), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4136 (
	.O(n3484),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_15__7_),
	.B1(n3500),
	.B2(Mfifo_xin_M_ffmem_mem_3__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4137 (
	.O(n3483),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_1__7_),
	.B1(n3502),
	.B2(Mfifo_xin_M_ffmem_mem_13__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4138 (
	.O(n3482),
	.A1(n3497),
	.A2(Mfifo_xin_M_ffmem_mem_7__7_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_5__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4139 (
	.O(n3481),
	.A1(n3495),
	.A2(Mfifo_xin_M_ffmem_mem_11__7_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_9__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4140 (
	.O(n3490),
	.I1(n3484),
	.I2(n3483),
	.I3(n3482),
	.I4(n3481), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4141 (
	.O(n3488),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_14__7_),
	.B1(n3497),
	.B2(Mfifo_xin_M_ffmem_mem_6__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4142 (
	.O(n3487),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_0__7_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_4__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4143 (
	.O(n3486),
	.A1(n3502),
	.A2(Mfifo_xin_M_ffmem_mem_12__7_),
	.B1(n3495),
	.B2(Mfifo_xin_M_ffmem_mem_10__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4144 (
	.O(n3485),
	.A1(n3500),
	.A2(Mfifo_xin_M_ffmem_mem_2__7_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_8__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4145 (
	.O(n3489),
	.I1(n3488),
	.I2(n3487),
	.I3(n3486),
	.I4(n3485), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4146 (
	.O(n2091),
	.A1(n3490),
	.A2(n3510),
	.B1(n3509),
	.B2(int_xin[7]),
	.C1(n3489),
	.C2(n3507), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4147 (
	.O(n3494),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_15__0_),
	.B1(n3495),
	.B2(Mfifo_xin_M_ffmem_mem_11__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4148 (
	.O(n3493),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_1__0_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_9__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4149 (
	.O(n3492),
	.A1(n3497),
	.A2(Mfifo_xin_M_ffmem_mem_7__0_),
	.B1(n3500),
	.B2(Mfifo_xin_M_ffmem_mem_3__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4150 (
	.O(n3491),
	.A1(n3502),
	.A2(Mfifo_xin_M_ffmem_mem_13__0_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_5__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4151 (
	.O(n3511),
	.I1(n3494),
	.I2(n3493),
	.I3(n3492),
	.I4(n3491), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4152 (
	.O(n3506),
	.A1(n3496),
	.A2(Mfifo_xin_M_ffmem_mem_0__0_),
	.B1(n3495),
	.B2(Mfifo_xin_M_ffmem_mem_10__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4153 (
	.O(n3505),
	.A1(n3498),
	.A2(Mfifo_xin_M_ffmem_mem_14__0_),
	.B1(n3497),
	.B2(Mfifo_xin_M_ffmem_mem_6__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4154 (
	.O(n3504),
	.A1(n3500),
	.A2(Mfifo_xin_M_ffmem_mem_2__0_),
	.B1(n3499),
	.B2(Mfifo_xin_M_ffmem_mem_4__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4155 (
	.O(n3503),
	.A1(n3502),
	.A2(Mfifo_xin_M_ffmem_mem_12__0_),
	.B1(n3501),
	.B2(Mfifo_xin_M_ffmem_mem_8__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4156 (
	.O(n3508),
	.I1(n3506),
	.I2(n3505),
	.I3(n3504),
	.I4(n3503), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO222X05AR9 U4157 (
	.O(n2090),
	.A1(n3511),
	.A2(n3510),
	.B1(n3509),
	.B2(int_xin[0]),
	.C1(n3508),
	.C2(n3507), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X05AR9 U4158 (
	.O(n3521),
	.B2(Mcntl_Mcntldata_c_W_r4[0]),
	.I1(n3512), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4159 (
	.O(n3517),
	.I(Mcntl_Mcntldata_c_W_r4[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12X05AR9 U4160 (
	.O(n3515),
	.A1(n3513),
	.B1(n3523),
	.B2(n3514), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI13X05AR9 U4161 (
	.O(n3516),
	.A1(n3522),
	.B1(Mcntl_Mcntldata_c_W_d4[1]),
	.B2(n3524),
	.B3(n3515), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4162 (
	.O(n2088),
	.A1(n3526),
	.B1(n3516),
	.C1(n3521),
	.C2(n3517), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AO12X05AR9 U4163 (
	.O(n2081),
	.A1(n3518),
	.B1(n3519),
	.B2(Mcntl_Mcntldata_c_x_cin[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4164 (
	.O(n3527),
	.A1(n3521),
	.A2(Mcntl_Mcntldata_c_W_r4[1]),
	.B1(Mcntl_Mcntldata_c_W_r4[0]),
	.B2(n3520), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI13X05AR9 U4165 (
	.O(n3525),
	.A1(n3522),
	.B1(Mcntl_Mcntldata_c_W_d4[1]),
	.B2(n3524),
	.B3(n3523), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND3X05AR9 U4166 (
	.O(n2080),
	.I1(n3527),
	.I2(n3526),
	.I3(n3525), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X05AR9 U4167 (
	.O(n3534),
	.I1(n3529),
	.I2(n3528), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4168 (
	.O(n3531),
	.I1(Mcntl_Mcntldata_count[0]),
	.I2(n3530), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI22X05AR9 U4169 (
	.O(n2079),
	.A1(n3534),
	.A2(n3533),
	.B1(n3532),
	.B2(n3531), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4170 (
	.O(n3551),
	.I(n3535), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4171 (
	.O(n3548),
	.I(Mfifo_psum_waddr[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   CLKNOR2X1AR9 U4172 (
	.O(n3812),
	.I1(n3551),
	.I2(n3546), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U4173 (
	.O(n3793),
	.I(n3812), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR3X05AR9 U4174 (
	.O(n3780),
	.I1(sel_reg[0]),
	.I2(n3537),
	.I3(n3622), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR3X05AR9 U4175 (
	.O(n3711),
	.I1(n3805),
	.I2(n3537),
	.I3(n3536), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX1AR9 U4176 (
	.O(n3802),
	.I(n3711), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4177 (
	.O(n3541),
	.A1(n3802),
	.A2(psum1_reg2[0]),
	.B1(n2407),
	.B2(psum2_reg4[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4178 (
	.O(n3540),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[0]),
	.C1(n3805),
	.C2(psum4_reg2[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1OAR9 U4179 (
	.O(n3803),
	.I1(sel_reg[1]),
	.I2(n3536), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4180 (
	.O(n3539),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[0]),
	.C1(n3805),
	.C2(psum3_reg2[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR3X1AR9 U4181 (
	.O(n3751),
	.I1(sel_ccp),
	.I2(n3537),
	.I3(n3536), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4182 (
	.O(n3538),
	.I1(n3751),
	.I2(psum1_reg4[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4183 (
	.O(n3542),
	.I1(n3541),
	.I2(n3540),
	.I3(n3539),
	.I4(n3538), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4184 (
	.O(n3557),
	.A1(n3542),
	.B1(n3811),
	.B2(psum2_reg2[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4185 (
	.O(n2065),
	.A1(n3793),
	.A2(n3557),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4186 (
	.O(n3545),
	.I1(n3550),
	.I2(n3543), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4187 (
	.O(n2064),
	.A1(n3813),
	.A2(n3557),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OR2B1X05AR9 U4188 (
	.O(n3552),
	.B2(Mfifo_psum_waddr[1]),
	.I1(Mfifo_psum_waddr[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1OAR9 U4189 (
	.O(n3815),
	.I1(n3546),
	.I2(n3552), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4190 (
	.O(n2063),
	.A1(n3814),
	.A2(n3557),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U4191 (
	.O(n3794),
	.I1(n3545),
	.I2(n3552), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4192 (
	.O(n2062),
	.A1(n3794),
	.A2(n3557),
	.B1B(n3794),
	.B2B(Mfifo_psum_M_ffmem_mem_3__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4193 (
	.O(n3554),
	.I1(Mfifo_psum_waddr[2]),
	.I2(n3544), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   CLKNOR2X1AR9 U4194 (
	.O(n3816),
	.I1(n3546),
	.I2(n3554), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U4195 (
	.O(n3795),
	.I(n3816), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4196 (
	.O(n2061),
	.A1(n3795),
	.A2(n3557),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4197 (
	.O(n2060),
	.A1(n3817),
	.A2(n3557),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NOR2X1AR9 U4198 (
	.O(n3818),
	.I1(n3556),
	.I2(n3546), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4199 (
	.O(n2059),
	.A1(n2399),
	.A2(n3557),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND2B1X1AR9 U4200 (
	.O(n3738),
	.B2(Mfifo_psum_waddr[3]),
	.I1(n3547), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX1AR9 U4201 (
	.O(n3819),
	.I(n3738), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4202 (
	.O(n2058),
	.A1(n3819),
	.A2(n3557),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4203 (
	.O(n2057),
	.A1(n2400),
	.A2(n3557),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4204 (
	.O(n3553),
	.I1(n3550),
	.I2(Mfifo_psum_waddr[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4205 (
	.O(n2056),
	.A1(n3821),
	.A2(n3557),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   CLKNOR2X1AR9 U4206 (
	.O(n3796),
	.I1(n3552),
	.I2(n3555), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U4207 (
	.O(n3822),
	.I(n3796), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4208 (
	.O(n2055),
	.A1(n3822),
	.A2(n3557),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4209 (
	.O(n2054),
	.A1(n3797),
	.A2(n3557),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   CLKNOR2X1AR9 U4210 (
	.O(n3823),
	.I1(n3554),
	.I2(n3555), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U4211 (
	.O(n3798),
	.I(n3823), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4212 (
	.O(n2053),
	.A1(n3798),
	.A2(n3557),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4213 (
	.O(n2052),
	.A1(n3799),
	.A2(n3557),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   CLKNOR2X1AR9 U4214 (
	.O(n3825),
	.I1(n3556),
	.I2(n3555), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4215 (
	.O(n2051),
	.A1(n3825),
	.A2(n3557),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__21_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4216 (
	.O(n2050),
	.A1(n3801),
	.A2(n3557),
	.B1B(Mfifo_psum_M_ffmem_mem_15__21_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4217 (
	.O(n3562),
	.A1(n3558),
	.A2(psum1_reg4[1]),
	.B1(n3802),
	.B2(psum1_reg2[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4218 (
	.O(n3561),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[1]),
	.C1(n3805),
	.C2(psum3_reg2[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4219 (
	.O(n3560),
	.I1(n2407),
	.I2(psum2_reg4[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4220 (
	.O(n3559),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[1]),
	.C1(n3805),
	.C2(psum4_reg2[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4221 (
	.O(n3563),
	.I1(n3562),
	.I2(n3561),
	.I3(n3560),
	.I4(n3559), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4222 (
	.O(n2049),
	.A1(n3812),
	.A2(n3564),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4223 (
	.O(n2048),
	.A1(n3813),
	.A2(n3564),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4224 (
	.O(n2047),
	.A1(n3815),
	.A2(n3564),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4225 (
	.O(n2046),
	.A1(n3794),
	.A2(n3564),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4226 (
	.O(n2045),
	.A1(n3816),
	.A2(n3564),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4227 (
	.O(n2044),
	.A1(n3817),
	.A2(n3564),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4228 (
	.O(n2043),
	.A1(n3818),
	.A2(n3564),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4229 (
	.O(n2042),
	.A1(n3738),
	.A2(n3564),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4230 (
	.O(n2041),
	.A1(n3820),
	.A2(n3564),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4231 (
	.O(n2040),
	.A1(n3821),
	.A2(n3564),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4232 (
	.O(n2039),
	.A1(n3796),
	.A2(n3564),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4233 (
	.O(n2038),
	.A1(n3797),
	.A2(n3564),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4234 (
	.O(n2037),
	.A1(n3823),
	.A2(n3564),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4235 (
	.O(n2036),
	.A1(n3799),
	.A2(n3564),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4236 (
	.O(n2035),
	.A1(n3825),
	.A2(n3564),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__22_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4237 (
	.O(n2034),
	.A1(n3801),
	.A2(n3564),
	.B1B(Mfifo_psum_M_ffmem_mem_15__22_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4238 (
	.O(n3568),
	.A1(n3558),
	.A2(psum1_reg4[2]),
	.B1(n2407),
	.B2(psum2_reg4[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4239 (
	.O(n3567),
	.A1(n3811),
	.A2(psum2_reg2[2]),
	.B1(n3802),
	.B2(psum1_reg2[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4240 (
	.O(n3566),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[2]),
	.C1(n3805),
	.C2(psum4_reg2[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4241 (
	.O(n3565),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[2]),
	.C1(n3805),
	.C2(psum3_reg2[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U4242 (
	.O(n3569),
	.I1(n3568),
	.I2(n3567),
	.I3(n3566),
	.I4(n3565), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4243 (
	.O(n2033),
	.A1(n3812),
	.A2(n3569),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4244 (
	.O(n2032),
	.A1(n3813),
	.A2(n3569),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX1AR9 U4245 (
	.O(n3814),
	.I(n3815), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4246 (
	.O(n2031),
	.A1(n3815),
	.A2(n3569),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4247 (
	.O(n2030),
	.A1(n3794),
	.A2(n3569),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4248 (
	.O(n2029),
	.A1(n3816),
	.A2(n3569),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4249 (
	.O(n2028),
	.A1(n3817),
	.A2(n3569),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4250 (
	.O(n2027),
	.A1(n3818),
	.A2(n3569),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4251 (
	.O(n2026),
	.A1(n3738),
	.A2(n3569),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4252 (
	.O(n2025),
	.A1(n3820),
	.A2(n3569),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4253 (
	.O(n2024),
	.A1(n3821),
	.A2(n3569),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4254 (
	.O(n2023),
	.A1(n3796),
	.A2(n3569),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4255 (
	.O(n2022),
	.A1(n3797),
	.A2(n3569),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4256 (
	.O(n2021),
	.A1(n3823),
	.A2(n3569),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4257 (
	.O(n2020),
	.A1(n3799),
	.A2(n3569),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   BUFX05AR9 U4258 (
	.O(n3824),
	.I(n3825), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4259 (
	.O(n2019),
	.A1(n3825),
	.A2(n3569),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__23_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4260 (
	.O(n2018),
	.A1(n3801),
	.A2(n3569),
	.B1B(Mfifo_psum_M_ffmem_mem_15__23_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4261 (
	.O(n3573),
	.A1(n3558),
	.A2(psum1_reg4[3]),
	.B1(n3802),
	.B2(psum1_reg2[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4262 (
	.O(n3572),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[3]),
	.C1(n3805),
	.C2(psum4_reg2[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4263 (
	.O(n3571),
	.I1(n3811),
	.I2(psum2_reg2[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4264 (
	.O(n3570),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[3]),
	.C1(n3805),
	.C2(psum3_reg2[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4265 (
	.O(n3574),
	.I1(n3573),
	.I2(n3572),
	.I3(n3571),
	.I4(n3570), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4266 (
	.O(n3575),
	.A1(n3574),
	.B1(n2407),
	.B2(psum2_reg4[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4267 (
	.O(n2017),
	.A1(n3812),
	.A2(n3575),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4268 (
	.O(n2016),
	.A1(n3813),
	.A2(n3575),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4269 (
	.O(n2015),
	.A1(n3814),
	.A2(n3575),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4270 (
	.O(n2014),
	.A1(n3794),
	.A2(n3575),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4271 (
	.O(n2013),
	.A1(n3816),
	.A2(n3575),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4272 (
	.O(n2012),
	.A1(n3817),
	.A2(n3575),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4273 (
	.O(n2011),
	.A1(n2399),
	.A2(n3575),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4274 (
	.O(n2010),
	.A1(n3819),
	.A2(n3575),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4275 (
	.O(n2009),
	.A1(n2400),
	.A2(n3575),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4276 (
	.O(n2008),
	.A1(n3821),
	.A2(n3575),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4277 (
	.O(n2007),
	.A1(n3822),
	.A2(n3575),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4278 (
	.O(n2006),
	.A1(n3797),
	.A2(n3575),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4279 (
	.O(n2005),
	.A1(n3823),
	.A2(n3575),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4280 (
	.O(n2004),
	.A1(n3799),
	.A2(n3575),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4281 (
	.O(n2003),
	.A1(n3824),
	.A2(n3575),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__24_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4282 (
	.O(n2002),
	.A1(n3801),
	.A2(n3575),
	.B1B(Mfifo_psum_M_ffmem_mem_15__24_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   LOWMUX2X05AR9 U4283 (
	.O(n3580),
	.EB(n3776),
	.I0(psum4_reg4[4]),
	.I1(psum4_reg2[4]),
	.S(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4284 (
	.O(n3578),
	.I(psum2_reg2[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4285 (
	.O(n3577),
	.A1(n3802),
	.A2(psum1_reg2[4]),
	.B1(n2407),
	.B2(psum2_reg4[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4286 (
	.O(n3576),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[4]),
	.C1(n3805),
	.C2(psum3_reg2[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4287 (
	.O(n3579),
	.A1(n3577),
	.B1(n3576),
	.C1(n3578),
	.C2(n3780), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4288 (
	.O(n2001),
	.A1(n3812),
	.A2(n3581),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4289 (
	.O(n2000),
	.A1(n3813),
	.A2(n3581),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4290 (
	.O(n1999),
	.A1(n3814),
	.A2(n3581),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4291 (
	.O(n1998),
	.A1(n3794),
	.A2(n3581),
	.B1B(n3794),
	.B2B(Mfifo_psum_M_ffmem_mem_3__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4292 (
	.O(n1997),
	.A1(n3816),
	.A2(n3581),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4293 (
	.O(n1996),
	.A1(n3817),
	.A2(n3581),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4294 (
	.O(n1995),
	.A1(n2399),
	.A2(n3581),
	.B1B(n3818),
	.B2B(Mfifo_psum_M_ffmem_mem_6__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4295 (
	.O(n1994),
	.A1(n3819),
	.A2(n3581),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4296 (
	.O(n1993),
	.A1(n2400),
	.A2(n3581),
	.B1B(n3820),
	.B2B(Mfifo_psum_M_ffmem_mem_8__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4297 (
	.O(n1992),
	.A1(n3821),
	.A2(n3581),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4298 (
	.O(n1991),
	.A1(n3796),
	.A2(n3581),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4299 (
	.O(n1990),
	.A1(n3797),
	.A2(n3581),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4300 (
	.O(n1989),
	.A1(n3823),
	.A2(n3581),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4301 (
	.O(n1988),
	.A1(n3799),
	.A2(n3581),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4302 (
	.O(n1987),
	.A1(n3824),
	.A2(n3581),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__25_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4303 (
	.O(n1986),
	.A1(n3801),
	.A2(n3581),
	.B1B(Mfifo_psum_M_ffmem_mem_15__25_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4304 (
	.O(n3585),
	.A1(n3558),
	.A2(psum1_reg4[5]),
	.B1(n2407),
	.B2(psum2_reg4[5]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4305 (
	.O(n3584),
	.A1(n3811),
	.A2(psum2_reg2[5]),
	.B1(n3802),
	.B2(psum1_reg2[5]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4306 (
	.O(n3622),
	.I(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4307 (
	.O(n3583),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[5]),
	.C1(n3622),
	.C2(psum4_reg2[5]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4308 (
	.O(n3582),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[5]),
	.C1(n3622),
	.C2(psum3_reg2[5]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U4309 (
	.O(n3586),
	.I1(n3585),
	.I2(n3584),
	.I3(n3583),
	.I4(n3582), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4310 (
	.O(n1985),
	.A1(n3793),
	.A2(n3586),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4311 (
	.O(n1984),
	.A1(n3813),
	.A2(n3586),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4312 (
	.O(n1983),
	.A1(n3814),
	.A2(n3586),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4313 (
	.O(n1982),
	.A1(n3794),
	.A2(n3586),
	.B1B(n3794),
	.B2B(Mfifo_psum_M_ffmem_mem_3__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4314 (
	.O(n1981),
	.A1(n3795),
	.A2(n3586),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4315 (
	.O(n1980),
	.A1(n3817),
	.A2(n3586),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4316 (
	.O(n1979),
	.A1(n2399),
	.A2(n3586),
	.B1B(n3818),
	.B2B(Mfifo_psum_M_ffmem_mem_6__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4317 (
	.O(n1978),
	.A1(n3819),
	.A2(n3586),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4318 (
	.O(n1977),
	.A1(n2400),
	.A2(n3586),
	.B1B(n3820),
	.B2B(Mfifo_psum_M_ffmem_mem_8__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4319 (
	.O(n1976),
	.A1(n3821),
	.A2(n3586),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4320 (
	.O(n1975),
	.A1(n3796),
	.A2(n3586),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4321 (
	.O(n1974),
	.A1(n3797),
	.A2(n3586),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4322 (
	.O(n1973),
	.A1(n3798),
	.A2(n3586),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4323 (
	.O(n1972),
	.A1(n3799),
	.A2(n3586),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4324 (
	.O(n1971),
	.A1(n3825),
	.A2(n3586),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__26_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4325 (
	.O(n1970),
	.A1(n3801),
	.A2(n3586),
	.B1B(Mfifo_psum_M_ffmem_mem_15__26_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4326 (
	.O(n3590),
	.A1(n3802),
	.A2(psum1_reg2[6]),
	.B1(n2407),
	.B2(psum2_reg4[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4327 (
	.O(n3589),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[6]),
	.C1(n3622),
	.C2(psum3_reg2[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4328 (
	.O(n3588),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[6]),
	.C1(n3622),
	.C2(psum4_reg2[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4329 (
	.O(n3587),
	.I1(n3751),
	.I2(psum1_reg4[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4330 (
	.O(n3591),
	.I1(n3590),
	.I2(n3589),
	.I3(n3588),
	.I4(n3587), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4331 (
	.O(n3592),
	.A1(n3591),
	.B1(n3811),
	.B2(psum2_reg2[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4332 (
	.O(n1969),
	.A1(n3793),
	.A2(n3592),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4333 (
	.O(n1968),
	.A1(n3813),
	.A2(n3592),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4334 (
	.O(n1967),
	.A1(n3814),
	.A2(n3592),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4335 (
	.O(n1966),
	.A1(n3794),
	.A2(n3592),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4336 (
	.O(n1965),
	.A1(n3795),
	.A2(n3592),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4337 (
	.O(n1964),
	.A1(n3817),
	.A2(n3592),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4338 (
	.O(n1963),
	.A1(n2399),
	.A2(n3592),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4339 (
	.O(n1962),
	.A1(n3819),
	.A2(n3592),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4340 (
	.O(n1961),
	.A1(n2400),
	.A2(n3592),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4341 (
	.O(n1960),
	.A1(n3821),
	.A2(n3592),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4342 (
	.O(n1959),
	.A1(n3796),
	.A2(n3592),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4343 (
	.O(n1958),
	.A1(n3797),
	.A2(n3592),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4344 (
	.O(n1957),
	.A1(n3798),
	.A2(n3592),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4345 (
	.O(n1956),
	.A1(n3799),
	.A2(n3592),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4346 (
	.O(n1955),
	.A1(n3825),
	.A2(n3592),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__27_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4347 (
	.O(n1954),
	.A1(n3801),
	.A2(n3592),
	.B1B(Mfifo_psum_M_ffmem_mem_15__27_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4348 (
	.O(n3596),
	.A1(n3802),
	.A2(psum1_reg2[7]),
	.B1(n2407),
	.B2(psum2_reg4[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4349 (
	.O(n3595),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[7]),
	.C1(n3622),
	.C2(psum3_reg2[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4350 (
	.O(n3594),
	.I1(n3811),
	.I2(psum2_reg2[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4351 (
	.O(n3593),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[7]),
	.C1(n3622),
	.C2(psum4_reg2[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4352 (
	.O(n3597),
	.I1(n3596),
	.I2(n3595),
	.I3(n3594),
	.I4(n3593), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4353 (
	.O(n3598),
	.A1(n3597),
	.B1(n3751),
	.B2(psum1_reg4[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4354 (
	.O(n1953),
	.A1(n3812),
	.A2(n3598),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4355 (
	.O(n1952),
	.A1(n3813),
	.A2(n3598),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4356 (
	.O(n1951),
	.A1(n3815),
	.A2(n3598),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4357 (
	.O(n1950),
	.A1(n3794),
	.A2(n3598),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4358 (
	.O(n1949),
	.A1(n3816),
	.A2(n3598),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4359 (
	.O(n1948),
	.A1(n3817),
	.A2(n3598),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4360 (
	.O(n1947),
	.A1(n3818),
	.A2(n3598),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4361 (
	.O(n1946),
	.A1(n3738),
	.A2(n3598),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4362 (
	.O(n1945),
	.A1(n3820),
	.A2(n3598),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4363 (
	.O(n1944),
	.A1(n3821),
	.A2(n3598),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4364 (
	.O(n1943),
	.A1(n3796),
	.A2(n3598),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4365 (
	.O(n1942),
	.A1(n3797),
	.A2(n3598),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4366 (
	.O(n1941),
	.A1(n3823),
	.A2(n3598),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4367 (
	.O(n1940),
	.A1(n3799),
	.A2(n3598),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4368 (
	.O(n1939),
	.A1(n3825),
	.A2(n3598),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__28_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4369 (
	.O(n1938),
	.A1(n3801),
	.A2(n3598),
	.B1B(Mfifo_psum_M_ffmem_mem_15__28_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4370 (
	.O(n3602),
	.A1(n3802),
	.A2(psum1_reg2[8]),
	.B1(n2407),
	.B2(psum2_reg4[8]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4371 (
	.O(n3601),
	.A1(n3811),
	.A2(psum2_reg2[8]),
	.B1(n3751),
	.B2(psum1_reg4[8]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4372 (
	.O(n3600),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[8]),
	.C1(n3622),
	.C2(psum3_reg2[8]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4373 (
	.O(n3599),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[8]),
	.C1(n3622),
	.C2(psum4_reg2[8]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U4374 (
	.O(n3603),
	.I1(n3602),
	.I2(n3601),
	.I3(n3600),
	.I4(n3599), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4375 (
	.O(n1937),
	.A1(n3812),
	.A2(n3603),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4376 (
	.O(n1936),
	.A1(n3813),
	.A2(n3603),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4377 (
	.O(n1935),
	.A1(n3815),
	.A2(n3603),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4378 (
	.O(n1934),
	.A1(n2398),
	.A2(n3603),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4379 (
	.O(n1933),
	.A1(n3816),
	.A2(n3603),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4380 (
	.O(n1932),
	.A1(n3817),
	.A2(n3603),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4381 (
	.O(n1931),
	.A1(n3818),
	.A2(n3603),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4382 (
	.O(n1930),
	.A1(n3819),
	.A2(n3603),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4383 (
	.O(n1929),
	.A1(n3820),
	.A2(n3603),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4384 (
	.O(n1928),
	.A1(n3821),
	.A2(n3603),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4385 (
	.O(n1927),
	.A1(n3796),
	.A2(n3603),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4386 (
	.O(n1926),
	.A1(n3797),
	.A2(n3603),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4387 (
	.O(n1925),
	.A1(n3823),
	.A2(n3603),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4388 (
	.O(n1924),
	.A1(n3799),
	.A2(n3603),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4389 (
	.O(n1923),
	.A1(n3825),
	.A2(n3603),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__29_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4390 (
	.O(n1922),
	.A1(n3801),
	.A2(n3603),
	.B1B(Mfifo_psum_M_ffmem_mem_15__29_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4391 (
	.O(n3607),
	.A1(n3811),
	.A2(psum2_reg2[9]),
	.B1(n2407),
	.B2(psum2_reg4[9]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4392 (
	.O(n3606),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[9]),
	.C1(n3622),
	.C2(psum4_reg2[9]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4393 (
	.O(n3605),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[9]),
	.C1(n3622),
	.C2(psum3_reg2[9]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4394 (
	.O(n3604),
	.I1(n3802),
	.I2(psum1_reg2[9]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4395 (
	.O(n3608),
	.I1(n3607),
	.I2(n3606),
	.I3(n3605),
	.I4(n3604), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4396 (
	.O(n3609),
	.A1(n3608),
	.B1(n3751),
	.B2(psum1_reg4[9]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4397 (
	.O(n1921),
	.A1(n3812),
	.A2(n3609),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4398 (
	.O(n1920),
	.A1(n3813),
	.A2(n3609),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4399 (
	.O(n1919),
	.A1(n3815),
	.A2(n3609),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4400 (
	.O(n1918),
	.A1(n2398),
	.A2(n3609),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4401 (
	.O(n1917),
	.A1(n3816),
	.A2(n3609),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4402 (
	.O(n1916),
	.A1(n3817),
	.A2(n3609),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4403 (
	.O(n1915),
	.A1(n3818),
	.A2(n3609),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4404 (
	.O(n1914),
	.A1(n3819),
	.A2(n3609),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4405 (
	.O(n1913),
	.A1(n3820),
	.A2(n3609),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4406 (
	.O(n1912),
	.A1(n3821),
	.A2(n3609),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4407 (
	.O(n1911),
	.A1(n3796),
	.A2(n3609),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4408 (
	.O(n1910),
	.A1(n3797),
	.A2(n3609),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4409 (
	.O(n1909),
	.A1(n3823),
	.A2(n3609),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4410 (
	.O(n1908),
	.A1(n3799),
	.A2(n3609),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4411 (
	.O(n1907),
	.A1(n3825),
	.A2(n3609),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__30_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4412 (
	.O(n1906),
	.A1(n3801),
	.A2(n3609),
	.B1B(Mfifo_psum_M_ffmem_mem_15__30_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4413 (
	.O(n3613),
	.A1(n3811),
	.A2(psum2_reg2[10]),
	.B1(n3751),
	.B2(psum1_reg4[10]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4414 (
	.O(n3612),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[10]),
	.C1(n3622),
	.C2(psum4_reg2[10]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4415 (
	.O(n3611),
	.I1(n2407),
	.I2(psum2_reg4[10]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4416 (
	.O(n3610),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[10]),
	.C1(n3622),
	.C2(psum3_reg2[10]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4417 (
	.O(n3614),
	.I1(n3613),
	.I2(n3612),
	.I3(n3611),
	.I4(n3610), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4418 (
	.O(n3615),
	.A1(n3614),
	.B1(n3802),
	.B2(psum1_reg2[10]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4419 (
	.O(n1905),
	.A1(n3812),
	.A2(n3615),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4420 (
	.O(n1904),
	.A1(n3813),
	.A2(n3615),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4421 (
	.O(n1903),
	.A1(n3814),
	.A2(n3615),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4422 (
	.O(n1902),
	.A1(n2398),
	.A2(n3615),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4423 (
	.O(n1901),
	.A1(n3816),
	.A2(n3615),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4424 (
	.O(n1900),
	.A1(n3817),
	.A2(n3615),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4425 (
	.O(n1899),
	.A1(n2399),
	.A2(n3615),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4426 (
	.O(n1898),
	.A1(n3819),
	.A2(n3615),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4427 (
	.O(n1897),
	.A1(n2400),
	.A2(n3615),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4428 (
	.O(n1896),
	.A1(n3821),
	.A2(n3615),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4429 (
	.O(n1895),
	.A1(n3796),
	.A2(n3615),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4430 (
	.O(n1894),
	.A1(n3797),
	.A2(n3615),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4431 (
	.O(n1893),
	.A1(n3823),
	.A2(n3615),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4432 (
	.O(n1892),
	.A1(n3799),
	.A2(n3615),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4433 (
	.O(n1891),
	.A1(n3824),
	.A2(n3615),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__31_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4434 (
	.O(n1890),
	.A1(n3801),
	.A2(n3615),
	.B1B(Mfifo_psum_M_ffmem_mem_15__31_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   LOWMUX2X05AR9 U4435 (
	.O(n3620),
	.EB(n3776),
	.I0(psum4_reg4[11]),
	.I1(psum4_reg2[11]),
	.S(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4436 (
	.O(n3618),
	.I(psum1_reg2[11]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4437 (
	.O(n3617),
	.A1(n3811),
	.A2(psum2_reg2[11]),
	.B1(n2407),
	.B2(psum2_reg4[11]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4438 (
	.O(n3616),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[11]),
	.C1(n3622),
	.C2(psum3_reg2[11]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4439 (
	.O(n3619),
	.A1(n3617),
	.B1(n3616),
	.C1(n3618),
	.C2(n3711), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4440 (
	.O(n1889),
	.A1(n3812),
	.A2(n3621),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4441 (
	.O(n1888),
	.A1(n3813),
	.A2(n3621),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4442 (
	.O(n1887),
	.A1(n3815),
	.A2(n3621),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4443 (
	.O(n1886),
	.A1(n2398),
	.A2(n3621),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4444 (
	.O(n1885),
	.A1(n3816),
	.A2(n3621),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4445 (
	.O(n1884),
	.A1(n3817),
	.A2(n3621),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4446 (
	.O(n1883),
	.A1(n3818),
	.A2(n3621),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4447 (
	.O(n1882),
	.A1(n3819),
	.A2(n3621),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4448 (
	.O(n1881),
	.A1(n3820),
	.A2(n3621),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4449 (
	.O(n1880),
	.A1(n3821),
	.A2(n3621),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4450 (
	.O(n1879),
	.A1(n3796),
	.A2(n3621),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4451 (
	.O(n1878),
	.A1(n3797),
	.A2(n3621),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4452 (
	.O(n1877),
	.A1(n3823),
	.A2(n3621),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4453 (
	.O(n1876),
	.A1(n3799),
	.A2(n3621),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4454 (
	.O(n1875),
	.A1(n3825),
	.A2(n3621),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__32_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4455 (
	.O(n1874),
	.A1(n3801),
	.A2(n3621),
	.B1B(Mfifo_psum_M_ffmem_mem_15__32_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4456 (
	.O(n3626),
	.A1(n3811),
	.A2(psum2_reg2[12]),
	.B1(n2407),
	.B2(psum2_reg4[12]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4457 (
	.O(n3625),
	.A1(n3558),
	.A2(psum1_reg4[12]),
	.B1(n3802),
	.B2(psum1_reg2[12]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4458 (
	.O(n3624),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[12]),
	.C1(n3622),
	.C2(psum3_reg2[12]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX1AR9 U4459 (
	.O(n3805),
	.I(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4460 (
	.O(n3623),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[12]),
	.C1(n3805),
	.C2(psum4_reg2[12]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U4461 (
	.O(n3627),
	.I1(n3626),
	.I2(n3625),
	.I3(n3624),
	.I4(n3623), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4462 (
	.O(n1873),
	.A1(n3812),
	.A2(n3627),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4463 (
	.O(n1872),
	.A1(n3813),
	.A2(n3627),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4464 (
	.O(n1871),
	.A1(n3815),
	.A2(n3627),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4465 (
	.O(n1870),
	.A1(n2398),
	.A2(n3627),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4466 (
	.O(n1869),
	.A1(n3816),
	.A2(n3627),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4467 (
	.O(n1868),
	.A1(n3817),
	.A2(n3627),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4468 (
	.O(n1867),
	.A1(n3818),
	.A2(n3627),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4469 (
	.O(n1866),
	.A1(n3738),
	.A2(n3627),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4470 (
	.O(n1865),
	.A1(n3820),
	.A2(n3627),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4471 (
	.O(n1864),
	.A1(n3821),
	.A2(n3627),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4472 (
	.O(n1863),
	.A1(n3796),
	.A2(n3627),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4473 (
	.O(n1862),
	.A1(n3797),
	.A2(n3627),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4474 (
	.O(n1861),
	.A1(n3823),
	.A2(n3627),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4475 (
	.O(n1860),
	.A1(n3799),
	.A2(n3627),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4476 (
	.O(n1859),
	.A1(n3825),
	.A2(n3627),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__33_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4477 (
	.O(n1858),
	.A1(n3801),
	.A2(n3627),
	.B1B(Mfifo_psum_M_ffmem_mem_15__33_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4478 (
	.O(n3631),
	.A1(n3802),
	.A2(psum1_reg2[13]),
	.B1(n2407),
	.B2(psum2_reg4[13]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4479 (
	.O(n3630),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[13]),
	.C1(n3805),
	.C2(psum4_reg2[13]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4480 (
	.O(n3629),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[13]),
	.C1(n3805),
	.C2(psum3_reg2[13]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4481 (
	.O(n3628),
	.I1(n3558),
	.I2(psum1_reg4[13]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4482 (
	.O(n3632),
	.I1(n3631),
	.I2(n3630),
	.I3(n3629),
	.I4(n3628), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4483 (
	.O(n3633),
	.A1(n3632),
	.B1(n3811),
	.B2(psum2_reg2[13]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4484 (
	.O(n1857),
	.A1(n3812),
	.A2(n3633),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4485 (
	.O(n1856),
	.A1(n3813),
	.A2(n3633),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4486 (
	.O(n1855),
	.A1(n3815),
	.A2(n3633),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4487 (
	.O(n1854),
	.A1(n2398),
	.A2(n3633),
	.B1B(n3794),
	.B2B(Mfifo_psum_M_ffmem_mem_3__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4488 (
	.O(n1853),
	.A1(n3816),
	.A2(n3633),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4489 (
	.O(n1852),
	.A1(n3817),
	.A2(n3633),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4490 (
	.O(n1851),
	.A1(n3818),
	.A2(n3633),
	.B1B(n3818),
	.B2B(Mfifo_psum_M_ffmem_mem_6__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4491 (
	.O(n1850),
	.A1(n3819),
	.A2(n3633),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4492 (
	.O(n1849),
	.A1(n3820),
	.A2(n3633),
	.B1B(n3820),
	.B2B(Mfifo_psum_M_ffmem_mem_8__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4493 (
	.O(n1848),
	.A1(n3821),
	.A2(n3633),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4494 (
	.O(n1847),
	.A1(n3796),
	.A2(n3633),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4495 (
	.O(n1846),
	.A1(n3797),
	.A2(n3633),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4496 (
	.O(n1845),
	.A1(n3823),
	.A2(n3633),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4497 (
	.O(n1844),
	.A1(n3799),
	.A2(n3633),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4498 (
	.O(n1843),
	.A1(n3825),
	.A2(n3633),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__34_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4499 (
	.O(n1842),
	.A1(n3801),
	.A2(n3633),
	.B1B(Mfifo_psum_M_ffmem_mem_15__34_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   LOWMUX2X05AR9 U4500 (
	.O(n3638),
	.EB(n3776),
	.I0(psum4_reg4[14]),
	.I1(psum4_reg2[14]),
	.S(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4501 (
	.O(n3636),
	.I(psum2_reg2[14]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4502 (
	.O(n3635),
	.A1(n3558),
	.A2(psum1_reg4[14]),
	.B1(n2407),
	.B2(psum2_reg4[14]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4503 (
	.O(n3634),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[14]),
	.C1(n3805),
	.C2(psum3_reg2[14]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4504 (
	.O(n3637),
	.A1(n3635),
	.B1(n3634),
	.C1(n3636),
	.C2(n3780), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4505 (
	.O(n1841),
	.A1(n3812),
	.A2(n3639),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4506 (
	.O(n1840),
	.A1(n3813),
	.A2(n3639),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4507 (
	.O(n1839),
	.A1(n3815),
	.A2(n3639),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4508 (
	.O(n1838),
	.A1(n2398),
	.A2(n3639),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4509 (
	.O(n1837),
	.A1(n3816),
	.A2(n3639),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4510 (
	.O(n1836),
	.A1(n3817),
	.A2(n3639),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4511 (
	.O(n1835),
	.A1(n3818),
	.A2(n3639),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4512 (
	.O(n1834),
	.A1(n3819),
	.A2(n3639),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4513 (
	.O(n1833),
	.A1(n3820),
	.A2(n3639),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4514 (
	.O(n1832),
	.A1(n3821),
	.A2(n3639),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4515 (
	.O(n1831),
	.A1(n3796),
	.A2(n3639),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4516 (
	.O(n1830),
	.A1(n3797),
	.A2(n3639),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4517 (
	.O(n1829),
	.A1(n3823),
	.A2(n3639),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4518 (
	.O(n1828),
	.A1(n3799),
	.A2(n3639),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4519 (
	.O(n1827),
	.A1(n3825),
	.A2(n3639),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__35_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4520 (
	.O(n1826),
	.A1(n3801),
	.A2(n3639),
	.B1B(Mfifo_psum_M_ffmem_mem_15__35_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA122X05AR9 U4521 (
	.O(n3645),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[15]),
	.C1(n3805),
	.C2(psum3_reg2[15]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4522 (
	.O(n3643),
	.I(psum2_reg2[15]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4523 (
	.O(n3642),
	.A1(n3802),
	.A2(psum1_reg2[15]),
	.B1(n2407),
	.B2(psum2_reg4[15]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4524 (
	.O(n3641),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[15]),
	.C1(n3805),
	.C2(psum4_reg2[15]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4525 (
	.O(n3644),
	.A1(n3642),
	.B1(n3641),
	.C1(n3780),
	.C2(n3643), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4526 (
	.O(n1825),
	.A1(n3812),
	.A2(n3646),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4527 (
	.O(n1824),
	.A1(n3813),
	.A2(n3646),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4528 (
	.O(n1823),
	.A1(n3815),
	.A2(n3646),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4529 (
	.O(n1822),
	.A1(n2398),
	.A2(n3646),
	.B1B(n3794),
	.B2B(Mfifo_psum_M_ffmem_mem_3__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4530 (
	.O(n1821),
	.A1(n3816),
	.A2(n3646),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4531 (
	.O(n1820),
	.A1(n3817),
	.A2(n3646),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4532 (
	.O(n1819),
	.A1(n3818),
	.A2(n3646),
	.B1B(n3818),
	.B2B(Mfifo_psum_M_ffmem_mem_6__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4533 (
	.O(n1818),
	.A1(n3819),
	.A2(n3646),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4534 (
	.O(n1817),
	.A1(n3820),
	.A2(n3646),
	.B1B(n3820),
	.B2B(Mfifo_psum_M_ffmem_mem_8__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4535 (
	.O(n1816),
	.A1(n3821),
	.A2(n3646),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4536 (
	.O(n1815),
	.A1(n3796),
	.A2(n3646),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4537 (
	.O(n1814),
	.A1(n3797),
	.A2(n3646),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4538 (
	.O(n1813),
	.A1(n3823),
	.A2(n3646),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4539 (
	.O(n1812),
	.A1(n3799),
	.A2(n3646),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4540 (
	.O(n1811),
	.A1(n3825),
	.A2(n3646),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__36_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4541 (
	.O(n1810),
	.A1(n3801),
	.A2(n3646),
	.B1B(Mfifo_psum_M_ffmem_mem_15__36_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4542 (
	.O(n3650),
	.A1(n3811),
	.A2(psum2_reg2[16]),
	.B1(n3558),
	.B2(psum1_reg4[16]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4543 (
	.O(n3649),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[16]),
	.C1(n3805),
	.C2(psum4_reg2[16]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4544 (
	.O(n3648),
	.I1(n3802),
	.I2(psum1_reg2[16]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4545 (
	.O(n3647),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[16]),
	.C1(n3805),
	.C2(psum3_reg2[16]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4546 (
	.O(n3651),
	.I1(n3650),
	.I2(n3649),
	.I3(n3648),
	.I4(n3647), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4547 (
	.O(n3652),
	.A1(n3651),
	.B1(n2407),
	.B2(psum2_reg4[16]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4548 (
	.O(n1809),
	.A1(n3812),
	.A2(n3652),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4549 (
	.O(n1808),
	.A1(n3813),
	.A2(n3652),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4550 (
	.O(n1807),
	.A1(n3815),
	.A2(n3652),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4551 (
	.O(n1806),
	.A1(n2398),
	.A2(n3652),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4552 (
	.O(n1805),
	.A1(n3816),
	.A2(n3652),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4553 (
	.O(n1804),
	.A1(n3817),
	.A2(n3652),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4554 (
	.O(n1803),
	.A1(n3818),
	.A2(n3652),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4555 (
	.O(n1802),
	.A1(n3738),
	.A2(n3652),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4556 (
	.O(n1801),
	.A1(n3820),
	.A2(n3652),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4557 (
	.O(n1800),
	.A1(n3821),
	.A2(n3652),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4558 (
	.O(n1799),
	.A1(n3796),
	.A2(n3652),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4559 (
	.O(n1798),
	.A1(n3797),
	.A2(n3652),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4560 (
	.O(n1797),
	.A1(n3823),
	.A2(n3652),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4561 (
	.O(n1796),
	.A1(n3799),
	.A2(n3652),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4562 (
	.O(n1795),
	.A1(n3825),
	.A2(n3652),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__37_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4563 (
	.O(n1794),
	.A1(n3801),
	.A2(n3652),
	.B1B(Mfifo_psum_M_ffmem_mem_15__37_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   LOWMUX2X05AR9 U4564 (
	.O(n3657),
	.EB(n3776),
	.I0(psum4_reg4[17]),
	.I1(psum4_reg2[17]),
	.S(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4565 (
	.O(n3655),
	.I(psum2_reg2[17]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4566 (
	.O(n3654),
	.A1(n3558),
	.A2(psum1_reg4[17]),
	.B1(n3802),
	.B2(psum1_reg2[17]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4567 (
	.O(n3653),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[17]),
	.C1(n3805),
	.C2(psum3_reg2[17]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4568 (
	.O(n3656),
	.A1(n3654),
	.B1(n3653),
	.C1(n3780),
	.C2(n3655), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4569 (
	.O(n1793),
	.A1(n3812),
	.A2(n3658),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4570 (
	.O(n1792),
	.A1(n3813),
	.A2(n3658),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4571 (
	.O(n1791),
	.A1(n3815),
	.A2(n3658),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4572 (
	.O(n1790),
	.A1(n2398),
	.A2(n3658),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4573 (
	.O(n1789),
	.A1(n3816),
	.A2(n3658),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4574 (
	.O(n1788),
	.A1(n3817),
	.A2(n3658),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4575 (
	.O(n1787),
	.A1(n3818),
	.A2(n3658),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4576 (
	.O(n1786),
	.A1(n3819),
	.A2(n3658),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4577 (
	.O(n1785),
	.A1(n3820),
	.A2(n3658),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4578 (
	.O(n1784),
	.A1(n3821),
	.A2(n3658),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4579 (
	.O(n1783),
	.A1(n3796),
	.A2(n3658),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4580 (
	.O(n1782),
	.A1(n3797),
	.A2(n3658),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4581 (
	.O(n1781),
	.A1(n3823),
	.A2(n3658),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4582 (
	.O(n1780),
	.A1(n3799),
	.A2(n3658),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4583 (
	.O(n1779),
	.A1(n3825),
	.A2(n3658),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__38_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4584 (
	.O(n1778),
	.A1(n3801),
	.A2(n3658),
	.B1B(Mfifo_psum_M_ffmem_mem_15__38_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4585 (
	.O(n3662),
	.A1(n3811),
	.A2(psum2_reg2[18]),
	.B1(n3802),
	.B2(psum1_reg2[18]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4586 (
	.O(n3661),
	.A1(n3558),
	.A2(psum1_reg4[18]),
	.B1(n2407),
	.B2(psum2_reg4[18]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4587 (
	.O(n3660),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[18]),
	.C1(n3805),
	.C2(psum4_reg2[18]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4588 (
	.O(n3659),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[18]),
	.C1(n3805),
	.C2(psum3_reg2[18]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U4589 (
	.O(n3663),
	.I1(n3662),
	.I2(n3661),
	.I3(n3660),
	.I4(n3659), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4590 (
	.O(n1777),
	.A1(n3812),
	.A2(n3663),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4591 (
	.O(n1776),
	.A1(n3813),
	.A2(n3663),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4592 (
	.O(n1775),
	.A1(n3815),
	.A2(n3663),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4593 (
	.O(n1774),
	.A1(n2398),
	.A2(n3663),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4594 (
	.O(n1773),
	.A1(n3816),
	.A2(n3663),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4595 (
	.O(n1772),
	.A1(n3817),
	.A2(n3663),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4596 (
	.O(n1771),
	.A1(n3818),
	.A2(n3663),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4597 (
	.O(n1770),
	.A1(n3738),
	.A2(n3663),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4598 (
	.O(n1769),
	.A1(n3820),
	.A2(n3663),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4599 (
	.O(n1768),
	.A1(n3821),
	.A2(n3663),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4600 (
	.O(n1767),
	.A1(n3796),
	.A2(n3663),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4601 (
	.O(n1766),
	.A1(n3797),
	.A2(n3663),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4602 (
	.O(n1765),
	.A1(n3823),
	.A2(n3663),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4603 (
	.O(n1764),
	.A1(n3799),
	.A2(n3663),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4604 (
	.O(n1763),
	.A1(n3825),
	.A2(n3663),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__39_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4605 (
	.O(n1762),
	.A1(n3801),
	.A2(n3663),
	.B1B(Mfifo_psum_M_ffmem_mem_15__39_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4606 (
	.O(n3667),
	.A1(n3558),
	.A2(psum1_reg4[19]),
	.B1(n3802),
	.B2(psum1_reg2[19]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4607 (
	.O(n3666),
	.A1(n3811),
	.A2(psum2_reg2[19]),
	.B1(n2407),
	.B2(psum2_reg4[19]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4608 (
	.O(n3665),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[19]),
	.C1(n3805),
	.C2(psum3_reg2[19]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4609 (
	.O(n3664),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[19]),
	.C1(n3805),
	.C2(psum4_reg2[19]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U4610 (
	.O(n3668),
	.I1(n3667),
	.I2(n3666),
	.I3(n3665),
	.I4(n3664), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4611 (
	.O(n1761),
	.A1(n3812),
	.A2(n3668),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4612 (
	.O(n1760),
	.A1(n3813),
	.A2(n3668),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4613 (
	.O(n1759),
	.A1(n3815),
	.A2(n3668),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4614 (
	.O(n1758),
	.A1(n2398),
	.A2(n3668),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4615 (
	.O(n1757),
	.A1(n3816),
	.A2(n3668),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4616 (
	.O(n1756),
	.A1(n3817),
	.A2(n3668),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4617 (
	.O(n1755),
	.A1(n3818),
	.A2(n3668),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4618 (
	.O(n1754),
	.A1(n3738),
	.A2(n3668),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4619 (
	.O(n1753),
	.A1(n3820),
	.A2(n3668),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4620 (
	.O(n1752),
	.A1(n3821),
	.A2(n3668),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4621 (
	.O(n1751),
	.A1(n3796),
	.A2(n3668),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4622 (
	.O(n1750),
	.A1(n3797),
	.A2(n3668),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4623 (
	.O(n1749),
	.A1(n3823),
	.A2(n3668),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4624 (
	.O(n1748),
	.A1(n3799),
	.A2(n3668),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4625 (
	.O(n1747),
	.A1(n3825),
	.A2(n3668),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__40_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4626 (
	.O(n1746),
	.A1(n3801),
	.A2(n3668),
	.B1B(Mfifo_psum_M_ffmem_mem_15__40_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4627 (
	.O(n3672),
	.A1(n3558),
	.A2(psum1_reg4[20]),
	.B1(n3802),
	.B2(psum1_reg2[20]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4628 (
	.O(n3671),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg4[20]),
	.C1(n3805),
	.C2(psum4_reg2[20]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4629 (
	.O(n3670),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg4[20]),
	.C1(n3805),
	.C2(psum3_reg2[20]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4630 (
	.O(n3669),
	.I1(n2407),
	.I2(psum2_reg4[20]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4631 (
	.O(n3673),
	.I1(n3672),
	.I2(n3671),
	.I3(n3670),
	.I4(n3669), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4632 (
	.O(n3674),
	.A1(n3673),
	.B1(n3811),
	.B2(psum2_reg2[20]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4633 (
	.O(n1745),
	.A1(n3812),
	.A2(n3674),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4634 (
	.O(n1744),
	.A1(n3813),
	.A2(n3674),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4635 (
	.O(n1743),
	.A1(n3815),
	.A2(n3674),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4636 (
	.O(n1742),
	.A1(n2398),
	.A2(n3674),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4637 (
	.O(n1741),
	.A1(n3816),
	.A2(n3674),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4638 (
	.O(n1740),
	.A1(n3817),
	.A2(n3674),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4639 (
	.O(n1739),
	.A1(n3818),
	.A2(n3674),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4640 (
	.O(n1738),
	.A1(n3819),
	.A2(n3674),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4641 (
	.O(n1737),
	.A1(n3820),
	.A2(n3674),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4642 (
	.O(n1736),
	.A1(n3821),
	.A2(n3674),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4643 (
	.O(n1735),
	.A1(n3796),
	.A2(n3674),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4644 (
	.O(n1734),
	.A1(n3797),
	.A2(n3674),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4645 (
	.O(n1733),
	.A1(n3823),
	.A2(n3674),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4646 (
	.O(n1732),
	.A1(n3799),
	.A2(n3674),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4647 (
	.O(n1731),
	.A1(n3825),
	.A2(n3674),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__41_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4648 (
	.O(n1730),
	.A1(n3801),
	.A2(n3674),
	.B1B(Mfifo_psum_M_ffmem_mem_15__41_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   LOWMUX2X05AR9 U4649 (
	.O(n3679),
	.EB(n3776),
	.I0(psum4_reg3[0]),
	.I1(psum4_reg1[0]),
	.S(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4650 (
	.O(n3677),
	.I(psum1_reg1[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4651 (
	.O(n3676),
	.A1(n3558),
	.A2(psum1_reg3[0]),
	.B1(n2407),
	.B2(psum2_reg3[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4652 (
	.O(n3675),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[0]),
	.C1(n3805),
	.C2(psum3_reg1[0]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4653 (
	.O(n3678),
	.A1(n3676),
	.B1(n3675),
	.C1(n3677),
	.C2(n3711), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4654 (
	.O(n1729),
	.A1(n3812),
	.A2(n3680),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4655 (
	.O(n1728),
	.A1(n3813),
	.A2(n3680),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4656 (
	.O(n1727),
	.A1(n3814),
	.A2(n3680),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4657 (
	.O(n1726),
	.A1(n2398),
	.A2(n3680),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4658 (
	.O(n1725),
	.A1(n3816),
	.A2(n3680),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4659 (
	.O(n1724),
	.A1(n3817),
	.A2(n3680),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4660 (
	.O(n1723),
	.A1(n2399),
	.A2(n3680),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4661 (
	.O(n1722),
	.A1(n3819),
	.A2(n3680),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4662 (
	.O(n1721),
	.A1(n2400),
	.A2(n3680),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4663 (
	.O(n1720),
	.A1(n3821),
	.A2(n3680),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4664 (
	.O(n1719),
	.A1(n3796),
	.A2(n3680),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4665 (
	.O(n1718),
	.A1(n3797),
	.A2(n3680),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4666 (
	.O(n1717),
	.A1(n3823),
	.A2(n3680),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4667 (
	.O(n1716),
	.A1(n3799),
	.A2(n3680),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4668 (
	.O(n1715),
	.A1(n3824),
	.A2(n3680),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__0_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4669 (
	.O(n1714),
	.A1(n3801),
	.A2(n3680),
	.B1B(Mfifo_psum_M_ffmem_mem_15__0_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4670 (
	.O(n3684),
	.A1(n3751),
	.A2(psum1_reg3[1]),
	.B1(n3802),
	.B2(psum1_reg1[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4671 (
	.O(n3683),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[1]),
	.C1(n3805),
	.C2(psum4_reg1[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4672 (
	.O(n3682),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[1]),
	.C1(psum3_reg1[1]),
	.C2(n3805), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4673 (
	.O(n3681),
	.I1(n2407),
	.I2(psum2_reg3[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4674 (
	.O(n3685),
	.I1(n3684),
	.I2(n3683),
	.I3(n3682),
	.I4(n3681), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4675 (
	.O(n1713),
	.A1(n3812),
	.A2(n3686),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4676 (
	.O(n1712),
	.A1(n3813),
	.A2(n3686),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4677 (
	.O(n1711),
	.A1(n3815),
	.A2(n3686),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4678 (
	.O(n1710),
	.A1(n2398),
	.A2(n3686),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4679 (
	.O(n1709),
	.A1(n3816),
	.A2(n3686),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4680 (
	.O(n1708),
	.A1(n3817),
	.A2(n3686),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4681 (
	.O(n1707),
	.A1(n3818),
	.A2(n3686),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4682 (
	.O(n1706),
	.A1(n3819),
	.A2(n3686),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4683 (
	.O(n1705),
	.A1(n3820),
	.A2(n3686),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4684 (
	.O(n1704),
	.A1(n3821),
	.A2(n3686),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4685 (
	.O(n1703),
	.A1(n3822),
	.A2(n3686),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4686 (
	.O(n1702),
	.A1(n3797),
	.A2(n3686),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4687 (
	.O(n1701),
	.A1(n3823),
	.A2(n3686),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4688 (
	.O(n1700),
	.A1(n3799),
	.A2(n3686),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4689 (
	.O(n1699),
	.A1(n3825),
	.A2(n3686),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__1_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4690 (
	.O(n1698),
	.A1(n3801),
	.A2(n3686),
	.B1B(Mfifo_psum_M_ffmem_mem_15__1_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4691 (
	.O(n3690),
	.A1(n3802),
	.A2(psum1_reg1[2]),
	.B1(n2407),
	.B2(psum2_reg3[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4692 (
	.O(n3689),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[2]),
	.C1(n3805),
	.C2(psum4_reg1[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4693 (
	.O(n3688),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[2]),
	.C1(n3805),
	.C2(psum3_reg1[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4694 (
	.O(n3687),
	.I1(n3811),
	.I2(psum2_reg1[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4695 (
	.O(n3691),
	.I1(n3690),
	.I2(n3689),
	.I3(n3688),
	.I4(n3687), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4696 (
	.O(n3692),
	.A1(n3691),
	.B1(n3751),
	.B2(psum1_reg3[2]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4697 (
	.O(n1697),
	.A1(n3812),
	.A2(n3692),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4698 (
	.O(n1696),
	.A1(n3813),
	.A2(n3692),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4699 (
	.O(n1695),
	.A1(n3814),
	.A2(n3692),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4700 (
	.O(n1694),
	.A1(n2398),
	.A2(n3692),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4701 (
	.O(n1693),
	.A1(n3816),
	.A2(n3692),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4702 (
	.O(n1692),
	.A1(n3817),
	.A2(n3692),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4703 (
	.O(n1691),
	.A1(n2399),
	.A2(n3692),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4704 (
	.O(n1690),
	.A1(n3819),
	.A2(n3692),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4705 (
	.O(n1689),
	.A1(n2400),
	.A2(n3692),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4706 (
	.O(n1688),
	.A1(n3821),
	.A2(n3692),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4707 (
	.O(n1687),
	.A1(n3822),
	.A2(n3692),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4708 (
	.O(n1686),
	.A1(n3797),
	.A2(n3692),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4709 (
	.O(n1685),
	.A1(n3823),
	.A2(n3692),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4710 (
	.O(n1684),
	.A1(n3799),
	.A2(n3692),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4711 (
	.O(n1683),
	.A1(n3824),
	.A2(n3692),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__2_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4712 (
	.O(n1682),
	.A1(n3801),
	.A2(n3692),
	.B1B(Mfifo_psum_M_ffmem_mem_15__2_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4713 (
	.O(n3696),
	.A1(n3811),
	.A2(psum2_reg1[3]),
	.B1(n3802),
	.B2(psum1_reg1[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4714 (
	.O(n3695),
	.A1(n3558),
	.A2(psum1_reg3[3]),
	.B1(n2407),
	.B2(psum2_reg3[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4715 (
	.O(n3694),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[3]),
	.C1(n3622),
	.C2(psum3_reg1[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4716 (
	.O(n3693),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[3]),
	.C1(n3622),
	.C2(psum4_reg1[3]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U4717 (
	.O(n3697),
	.I1(n3696),
	.I2(n3695),
	.I3(n3694),
	.I4(n3693), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4718 (
	.O(n1681),
	.A1(n3812),
	.A2(n3697),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4719 (
	.O(n1680),
	.A1(n3813),
	.A2(n3697),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4720 (
	.O(n1679),
	.A1(n3814),
	.A2(n3697),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4721 (
	.O(n1678),
	.A1(n2398),
	.A2(n3697),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4722 (
	.O(n1677),
	.A1(n3816),
	.A2(n3697),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4723 (
	.O(n1676),
	.A1(n3817),
	.A2(n3697),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4724 (
	.O(n1675),
	.A1(n2399),
	.A2(n3697),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4725 (
	.O(n1674),
	.A1(n3819),
	.A2(n3697),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4726 (
	.O(n1673),
	.A1(n2400),
	.A2(n3697),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4727 (
	.O(n1672),
	.A1(n3821),
	.A2(n3697),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4728 (
	.O(n1671),
	.A1(n3822),
	.A2(n3697),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4729 (
	.O(n1670),
	.A1(n3797),
	.A2(n3697),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4730 (
	.O(n1669),
	.A1(n3823),
	.A2(n3697),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4731 (
	.O(n1668),
	.A1(n3799),
	.A2(n3697),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4732 (
	.O(n1667),
	.A1(n3824),
	.A2(n3697),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__3_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4733 (
	.O(n1666),
	.A1(n3801),
	.A2(n3697),
	.B1B(Mfifo_psum_M_ffmem_mem_15__3_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4734 (
	.O(n3701),
	.A1(n3811),
	.A2(psum2_reg1[4]),
	.B1(n2407),
	.B2(psum2_reg3[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4735 (
	.O(n3700),
	.A1(n3751),
	.A2(psum1_reg3[4]),
	.B1(n3802),
	.B2(psum1_reg1[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4736 (
	.O(n3699),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[4]),
	.C1(n3622),
	.C2(psum4_reg1[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4737 (
	.O(n3698),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[4]),
	.C1(n3622),
	.C2(psum3_reg1[4]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U4738 (
	.O(n3702),
	.I1(n3701),
	.I2(n3700),
	.I3(n3699),
	.I4(n3698), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4739 (
	.O(n1665),
	.A1(n3793),
	.A2(n3702),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4740 (
	.O(n1664),
	.A1(n3813),
	.A2(n3702),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4741 (
	.O(n1663),
	.A1(n3814),
	.A2(n3702),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4742 (
	.O(n1662),
	.A1(n3794),
	.A2(n3702),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4743 (
	.O(n1661),
	.A1(n3795),
	.A2(n3702),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4744 (
	.O(n1660),
	.A1(n3817),
	.A2(n3702),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4745 (
	.O(n1659),
	.A1(n2399),
	.A2(n3702),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4746 (
	.O(n1658),
	.A1(n3819),
	.A2(n3702),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4747 (
	.O(n1657),
	.A1(n2400),
	.A2(n3702),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4748 (
	.O(n1656),
	.A1(n3821),
	.A2(n3702),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4749 (
	.O(n1655),
	.A1(n3822),
	.A2(n3702),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4750 (
	.O(n1654),
	.A1(n3797),
	.A2(n3702),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4751 (
	.O(n1653),
	.A1(n3798),
	.A2(n3702),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4752 (
	.O(n1652),
	.A1(n3799),
	.A2(n3702),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4753 (
	.O(n1651),
	.A1(n3825),
	.A2(n3702),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__4_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4754 (
	.O(n1650),
	.A1(n3801),
	.A2(n3702),
	.B1B(Mfifo_psum_M_ffmem_mem_15__4_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   LOWMUX2X05AR9 U4755 (
	.O(n3707),
	.EB(n3776),
	.I0(psum4_reg3[5]),
	.I1(psum4_reg1[5]),
	.S(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4756 (
	.O(n3705),
	.I(psum2_reg1[5]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4757 (
	.O(n3704),
	.A1(n3751),
	.A2(psum1_reg3[5]),
	.B1(n2407),
	.B2(psum2_reg3[5]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4758 (
	.O(n3703),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[5]),
	.C1(n3805),
	.C2(psum3_reg1[5]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4759 (
	.O(n3706),
	.A1(n3704),
	.B1(n3703),
	.C1(n3705),
	.C2(n3780), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U4760 (
	.O(n3708),
	.A1(n3707),
	.B1(n3706),
	.C1(n3802),
	.C2(psum1_reg1[5]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4761 (
	.O(n1649),
	.A1(n3793),
	.A2(n3708),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4762 (
	.O(n1648),
	.A1(n3813),
	.A2(n3708),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4763 (
	.O(n1647),
	.A1(n3814),
	.A2(n3708),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4764 (
	.O(n1646),
	.A1(n3794),
	.A2(n3708),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4765 (
	.O(n1645),
	.A1(n3795),
	.A2(n3708),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4766 (
	.O(n1644),
	.A1(n3817),
	.A2(n3708),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4767 (
	.O(n1643),
	.A1(n2399),
	.A2(n3708),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4768 (
	.O(n1642),
	.A1(n3819),
	.A2(n3708),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4769 (
	.O(n1641),
	.A1(n2400),
	.A2(n3708),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4770 (
	.O(n1640),
	.A1(n3821),
	.A2(n3708),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4771 (
	.O(n1639),
	.A1(n3822),
	.A2(n3708),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4772 (
	.O(n1638),
	.A1(n3797),
	.A2(n3708),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4773 (
	.O(n1637),
	.A1(n3798),
	.A2(n3708),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4774 (
	.O(n1636),
	.A1(n3799),
	.A2(n3708),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4775 (
	.O(n1635),
	.A1(n3825),
	.A2(n3708),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__5_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4776 (
	.O(n1634),
	.A1(n3801),
	.A2(n3708),
	.B1B(Mfifo_psum_M_ffmem_mem_15__5_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OA122X05AR9 U4777 (
	.O(n3714),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[6]),
	.C1(n3805),
	.C2(psum3_reg1[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4778 (
	.O(n3712),
	.I(psum1_reg1[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4779 (
	.O(n3710),
	.A1(n3811),
	.A2(psum2_reg1[6]),
	.B1(n2407),
	.B2(psum2_reg3[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4780 (
	.O(n3709),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[6]),
	.C1(n3805),
	.C2(psum4_reg1[6]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4781 (
	.O(n3713),
	.A1(n3710),
	.B1(n3709),
	.C1(n3712),
	.C2(n3711), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4782 (
	.O(n1633),
	.A1(n3793),
	.A2(n3715),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4783 (
	.O(n1632),
	.A1(n3813),
	.A2(n3715),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4784 (
	.O(n1631),
	.A1(n3814),
	.A2(n3715),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4785 (
	.O(n1630),
	.A1(n2398),
	.A2(n3715),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4786 (
	.O(n1629),
	.A1(n3795),
	.A2(n3715),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4787 (
	.O(n1628),
	.A1(n3817),
	.A2(n3715),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4788 (
	.O(n1627),
	.A1(n2399),
	.A2(n3715),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4789 (
	.O(n1626),
	.A1(n3819),
	.A2(n3715),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4790 (
	.O(n1625),
	.A1(n2400),
	.A2(n3715),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4791 (
	.O(n1624),
	.A1(n3821),
	.A2(n3715),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4792 (
	.O(n1623),
	.A1(n3822),
	.A2(n3715),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4793 (
	.O(n1622),
	.A1(n3797),
	.A2(n3715),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4794 (
	.O(n1621),
	.A1(n3798),
	.A2(n3715),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4795 (
	.O(n1620),
	.A1(n3799),
	.A2(n3715),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4796 (
	.O(n1619),
	.A1(n3825),
	.A2(n3715),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__6_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4797 (
	.O(n1618),
	.A1(n3801),
	.A2(n3715),
	.B1B(Mfifo_psum_M_ffmem_mem_15__6_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4798 (
	.O(n3719),
	.A1(n3811),
	.A2(psum2_reg1[7]),
	.B1(n3558),
	.B2(psum1_reg3[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4799 (
	.O(n3718),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[7]),
	.C1(n3805),
	.C2(psum3_reg1[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4800 (
	.O(n3717),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[7]),
	.C1(n3805),
	.C2(psum4_reg1[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4801 (
	.O(n3716),
	.I1(n2407),
	.I2(psum2_reg3[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4802 (
	.O(n3720),
	.I1(n3719),
	.I2(n3718),
	.I3(n3717),
	.I4(n3716), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4803 (
	.O(n3721),
	.A1(n3720),
	.B1(n3802),
	.B2(psum1_reg1[7]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4804 (
	.O(n1617),
	.A1(n3793),
	.A2(n3721),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4805 (
	.O(n1616),
	.A1(n3813),
	.A2(n3721),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4806 (
	.O(n1615),
	.A1(n3814),
	.A2(n3721),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4807 (
	.O(n1614),
	.A1(n2398),
	.A2(n3721),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4808 (
	.O(n1613),
	.A1(n3795),
	.A2(n3721),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4809 (
	.O(n1612),
	.A1(n3817),
	.A2(n3721),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4810 (
	.O(n1611),
	.A1(n2399),
	.A2(n3721),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4811 (
	.O(n1610),
	.A1(n3819),
	.A2(n3721),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4812 (
	.O(n1609),
	.A1(n2400),
	.A2(n3721),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4813 (
	.O(n1608),
	.A1(n3821),
	.A2(n3721),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4814 (
	.O(n1607),
	.A1(n3822),
	.A2(n3721),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4815 (
	.O(n1606),
	.A1(n3797),
	.A2(n3721),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4816 (
	.O(n1605),
	.A1(n3798),
	.A2(n3721),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4817 (
	.O(n1604),
	.A1(n3799),
	.A2(n3721),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4818 (
	.O(n1603),
	.A1(n3825),
	.A2(n3721),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__7_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4819 (
	.O(n1602),
	.A1(n3801),
	.A2(n3721),
	.B1B(Mfifo_psum_M_ffmem_mem_15__7_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   LOWMUX2X05AR9 U4820 (
	.O(n3726),
	.EB(n3776),
	.I0(psum4_reg3[8]),
	.I1(psum4_reg1[8]),
	.S(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4821 (
	.O(n3724),
	.I(psum2_reg1[8]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4822 (
	.O(n3723),
	.A1(n3802),
	.A2(psum1_reg1[8]),
	.B1(n2407),
	.B2(psum2_reg3[8]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4823 (
	.O(n3722),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[8]),
	.C1(n3805),
	.C2(psum3_reg1[8]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4824 (
	.O(n3725),
	.A1(n3723),
	.B1(n3722),
	.C1(n3780),
	.C2(n3724), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4825 (
	.O(n1601),
	.A1(n3793),
	.A2(n3727),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4826 (
	.O(n1600),
	.A1(n3813),
	.A2(n3727),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4827 (
	.O(n1599),
	.A1(n3814),
	.A2(n3727),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4828 (
	.O(n1598),
	.A1(n2398),
	.A2(n3727),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4829 (
	.O(n1597),
	.A1(n3795),
	.A2(n3727),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4830 (
	.O(n1596),
	.A1(n3817),
	.A2(n3727),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4831 (
	.O(n1595),
	.A1(n2399),
	.A2(n3727),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4832 (
	.O(n1594),
	.A1(n3819),
	.A2(n3727),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4833 (
	.O(n1593),
	.A1(n2400),
	.A2(n3727),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4834 (
	.O(n1592),
	.A1(n3821),
	.A2(n3727),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4835 (
	.O(n1591),
	.A1(n3822),
	.A2(n3727),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4836 (
	.O(n1590),
	.A1(n3797),
	.A2(n3727),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4837 (
	.O(n1589),
	.A1(n3798),
	.A2(n3727),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4838 (
	.O(n1588),
	.A1(n3799),
	.A2(n3727),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4839 (
	.O(n1587),
	.A1(n3825),
	.A2(n3727),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__8_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4840 (
	.O(n1586),
	.A1(n3801),
	.A2(n3727),
	.B1B(Mfifo_psum_M_ffmem_mem_15__8_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   LOWMUX2X05AR9 U4841 (
	.O(n3732),
	.EB(n3776),
	.I0(psum4_reg3[9]),
	.I1(psum4_reg1[9]),
	.S(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4842 (
	.O(n3730),
	.I(psum2_reg1[9]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4843 (
	.O(n3729),
	.A1(n3751),
	.A2(psum1_reg3[9]),
	.B1(n3802),
	.B2(psum1_reg1[9]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4844 (
	.O(n3728),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[9]),
	.C1(n3805),
	.C2(psum3_reg1[9]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4845 (
	.O(n3731),
	.A1(n3729),
	.B1(n3728),
	.C1(n3730),
	.C2(n3780), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4846 (
	.O(n1585),
	.A1(n3812),
	.A2(n3733),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4847 (
	.O(n1584),
	.A1(n3813),
	.A2(n3733),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4848 (
	.O(n1583),
	.A1(n3814),
	.A2(n3733),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4849 (
	.O(n1582),
	.A1(n3794),
	.A2(n3733),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4850 (
	.O(n1581),
	.A1(n3816),
	.A2(n3733),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4851 (
	.O(n1580),
	.A1(n3817),
	.A2(n3733),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4852 (
	.O(n1579),
	.A1(n2399),
	.A2(n3733),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4853 (
	.O(n1578),
	.A1(n3819),
	.A2(n3733),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4854 (
	.O(n1577),
	.A1(n2400),
	.A2(n3733),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4855 (
	.O(n1576),
	.A1(n3821),
	.A2(n3733),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4856 (
	.O(n1575),
	.A1(n3822),
	.A2(n3733),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4857 (
	.O(n1574),
	.A1(n3797),
	.A2(n3733),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4858 (
	.O(n1573),
	.A1(n3823),
	.A2(n3733),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4859 (
	.O(n1572),
	.A1(n3799),
	.A2(n3733),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4860 (
	.O(n1571),
	.A1(n3824),
	.A2(n3733),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__9_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4861 (
	.O(n1570),
	.A1(n3801),
	.A2(n3733),
	.B1B(Mfifo_psum_M_ffmem_mem_15__9_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4862 (
	.O(n3737),
	.A1(n3811),
	.A2(psum2_reg1[10]),
	.B1(n2407),
	.B2(psum2_reg3[10]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4863 (
	.O(n3736),
	.A1(n3751),
	.A2(psum1_reg3[10]),
	.B1(n3802),
	.B2(psum1_reg1[10]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4864 (
	.O(n3735),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[10]),
	.C1(n3805),
	.C2(psum4_reg1[10]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4865 (
	.O(n3734),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[10]),
	.C1(n3805),
	.C2(psum3_reg1[10]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U4866 (
	.O(n3739),
	.I1(n3737),
	.I2(n3736),
	.I3(n3735),
	.I4(n3734), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4867 (
	.O(n1569),
	.A1(n3812),
	.A2(n3739),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4868 (
	.O(n1568),
	.A1(n3813),
	.A2(n3739),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4869 (
	.O(n1567),
	.A1(n3815),
	.A2(n3739),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4870 (
	.O(n1566),
	.A1(n3794),
	.A2(n3739),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4871 (
	.O(n1565),
	.A1(n3816),
	.A2(n3739),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4872 (
	.O(n1564),
	.A1(n3817),
	.A2(n3739),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4873 (
	.O(n1563),
	.A1(n3818),
	.A2(n3739),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4874 (
	.O(n1562),
	.A1(n3738),
	.A2(n3739),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4875 (
	.O(n1561),
	.A1(n3820),
	.A2(n3739),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4876 (
	.O(n1560),
	.A1(n3821),
	.A2(n3739),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4877 (
	.O(n1559),
	.A1(n3822),
	.A2(n3739),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4878 (
	.O(n1558),
	.A1(n3797),
	.A2(n3739),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4879 (
	.O(n1557),
	.A1(n3823),
	.A2(n3739),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4880 (
	.O(n1556),
	.A1(n3799),
	.A2(n3739),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4881 (
	.O(n1555),
	.A1(n3825),
	.A2(n3739),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__10_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4882 (
	.O(n1554),
	.A1(n3801),
	.A2(n3739),
	.B1B(Mfifo_psum_M_ffmem_mem_15__10_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   LOWMUX2X05AR9 U4883 (
	.O(n3744),
	.EB(n3776),
	.I0(psum4_reg3[11]),
	.I1(psum4_reg1[11]),
	.S(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4884 (
	.O(n3742),
	.I(psum2_reg1[11]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4885 (
	.O(n3741),
	.A1(n3802),
	.A2(psum1_reg1[11]),
	.B1(n2407),
	.B2(psum2_reg3[11]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4886 (
	.O(n3740),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[11]),
	.C1(n3805),
	.C2(psum3_reg1[11]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4887 (
	.O(n3743),
	.A1(n3741),
	.B1(n3740),
	.C1(n3742),
	.C2(n3780), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U4888 (
	.O(n3745),
	.A1(n3744),
	.B1(n3743),
	.C1(n3751),
	.C2(psum1_reg3[11]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4889 (
	.O(n1553),
	.A1(n3812),
	.A2(n3745),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4890 (
	.O(n1552),
	.A1(n3813),
	.A2(n3745),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4891 (
	.O(n1551),
	.A1(n3814),
	.A2(n3745),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4892 (
	.O(n1550),
	.A1(n2398),
	.A2(n3745),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4893 (
	.O(n1549),
	.A1(n3816),
	.A2(n3745),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4894 (
	.O(n1548),
	.A1(n3817),
	.A2(n3745),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4895 (
	.O(n1547),
	.A1(n2399),
	.A2(n3745),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4896 (
	.O(n1546),
	.A1(n3819),
	.A2(n3745),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4897 (
	.O(n1545),
	.A1(n2400),
	.A2(n3745),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4898 (
	.O(n1544),
	.A1(n3821),
	.A2(n3745),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4899 (
	.O(n1543),
	.A1(n3822),
	.A2(n3745),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4900 (
	.O(n1542),
	.A1(n3797),
	.A2(n3745),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4901 (
	.O(n1541),
	.A1(n3823),
	.A2(n3745),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4902 (
	.O(n1540),
	.A1(n3799),
	.A2(n3745),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4903 (
	.O(n1539),
	.A1(n3824),
	.A2(n3745),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__11_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4904 (
	.O(n1538),
	.A1(n3801),
	.A2(n3745),
	.B1B(Mfifo_psum_M_ffmem_mem_15__11_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4905 (
	.O(n3749),
	.A1(n3811),
	.A2(psum2_reg1[12]),
	.B1(n2407),
	.B2(psum2_reg3[12]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4906 (
	.O(n3748),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[12]),
	.C1(n3805),
	.C2(psum3_reg1[12]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4907 (
	.O(n3747),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[12]),
	.C1(n3805),
	.C2(psum4_reg1[12]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4908 (
	.O(n3746),
	.I1(n3802),
	.I2(psum1_reg1[12]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4909 (
	.O(n3750),
	.I1(n3749),
	.I2(n3748),
	.I3(n3747),
	.I4(n3746), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4910 (
	.O(n3752),
	.A1(n3750),
	.B1(n3751),
	.B2(psum1_reg3[12]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4911 (
	.O(n1537),
	.A1(n3793),
	.A2(n3752),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4912 (
	.O(n1536),
	.A1(n3813),
	.A2(n3752),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4913 (
	.O(n1535),
	.A1(n3814),
	.A2(n3752),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4914 (
	.O(n1534),
	.A1(n3794),
	.A2(n3752),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4915 (
	.O(n1533),
	.A1(n3795),
	.A2(n3752),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4916 (
	.O(n1532),
	.A1(n3817),
	.A2(n3752),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4917 (
	.O(n1531),
	.A1(n2399),
	.A2(n3752),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4918 (
	.O(n1530),
	.A1(n3819),
	.A2(n3752),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4919 (
	.O(n1529),
	.A1(n2400),
	.A2(n3752),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4920 (
	.O(n1528),
	.A1(n3821),
	.A2(n3752),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4921 (
	.O(n1527),
	.A1(n3822),
	.A2(n3752),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4922 (
	.O(n1526),
	.A1(n3797),
	.A2(n3752),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4923 (
	.O(n1525),
	.A1(n3798),
	.A2(n3752),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4924 (
	.O(n1524),
	.A1(n3799),
	.A2(n3752),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4925 (
	.O(n1523),
	.A1(n3825),
	.A2(n3752),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__12_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4926 (
	.O(n1522),
	.A1(n3801),
	.A2(n3752),
	.B1B(Mfifo_psum_M_ffmem_mem_15__12_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4927 (
	.O(n3756),
	.A1(n3811),
	.A2(psum2_reg1[13]),
	.B1(n2407),
	.B2(psum2_reg3[13]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4928 (
	.O(n3755),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[13]),
	.C1(n3805),
	.C2(psum3_reg1[13]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4929 (
	.O(n3754),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[13]),
	.C1(n3805),
	.C2(psum4_reg1[13]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4930 (
	.O(n3753),
	.I1(n3558),
	.I2(psum1_reg3[13]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4931 (
	.O(n3757),
	.I1(n3756),
	.I2(n3755),
	.I3(n3754),
	.I4(n3753), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4932 (
	.O(n3758),
	.A1(n3757),
	.B1(n3802),
	.B2(psum1_reg1[13]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4933 (
	.O(n1521),
	.A1(n3793),
	.A2(n3758),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4934 (
	.O(n1520),
	.A1(n3813),
	.A2(n3758),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4935 (
	.O(n1519),
	.A1(n3814),
	.A2(n3758),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4936 (
	.O(n1518),
	.A1(n3794),
	.A2(n3758),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4937 (
	.O(n1517),
	.A1(n3795),
	.A2(n3758),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4938 (
	.O(n1516),
	.A1(n3817),
	.A2(n3758),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4939 (
	.O(n1515),
	.A1(n2399),
	.A2(n3758),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4940 (
	.O(n1514),
	.A1(n3819),
	.A2(n3758),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4941 (
	.O(n1513),
	.A1(n2400),
	.A2(n3758),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4942 (
	.O(n1512),
	.A1(n3821),
	.A2(n3758),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4943 (
	.O(n1511),
	.A1(n3822),
	.A2(n3758),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4944 (
	.O(n1510),
	.A1(n3797),
	.A2(n3758),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4945 (
	.O(n1509),
	.A1(n3798),
	.A2(n3758),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4946 (
	.O(n1508),
	.A1(n3799),
	.A2(n3758),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4947 (
	.O(n1507),
	.A1(n3825),
	.A2(n3758),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__13_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4948 (
	.O(n1506),
	.A1(n3801),
	.A2(n3758),
	.B1B(Mfifo_psum_M_ffmem_mem_15__13_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   LOWMUX2X05AR9 U4949 (
	.O(n3763),
	.EB(n3776),
	.I0(psum4_reg3[14]),
	.I1(psum4_reg1[14]),
	.S(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U4950 (
	.O(n3761),
	.I(psum2_reg1[14]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4951 (
	.O(n3760),
	.A1(n3751),
	.A2(psum1_reg3[14]),
	.B1(n2407),
	.B2(psum2_reg3[14]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4952 (
	.O(n3759),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[14]),
	.C1(n3805),
	.C2(psum3_reg1[14]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U4953 (
	.O(n3762),
	.A1(n3760),
	.B1(n3759),
	.C1(n3780),
	.C2(n3761), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI112X05AR9 U4954 (
	.O(n3764),
	.A1(n3763),
	.B1(n3762),
	.C1(psum1_reg1[14]),
	.C2(n3802), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4955 (
	.O(n1505),
	.A1(n3812),
	.A2(n3764),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4956 (
	.O(n1504),
	.A1(n3813),
	.A2(n3764),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4957 (
	.O(n1503),
	.A1(n3815),
	.A2(n3764),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4958 (
	.O(n1502),
	.A1(n2398),
	.A2(n3764),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4959 (
	.O(n1501),
	.A1(n3816),
	.A2(n3764),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4960 (
	.O(n1500),
	.A1(n3817),
	.A2(n3764),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4961 (
	.O(n1499),
	.A1(n3818),
	.A2(n3764),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4962 (
	.O(n1498),
	.A1(n3819),
	.A2(n3764),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4963 (
	.O(n1497),
	.A1(n3820),
	.A2(n3764),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4964 (
	.O(n1496),
	.A1(n3821),
	.A2(n3764),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4965 (
	.O(n1495),
	.A1(n3822),
	.A2(n3764),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4966 (
	.O(n1494),
	.A1(n3797),
	.A2(n3764),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4967 (
	.O(n1493),
	.A1(n3823),
	.A2(n3764),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4968 (
	.O(n1492),
	.A1(n3799),
	.A2(n3764),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4969 (
	.O(n1491),
	.A1(n3825),
	.A2(n3764),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__14_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4970 (
	.O(n1490),
	.A1(n3801),
	.A2(n3764),
	.B1B(Mfifo_psum_M_ffmem_mem_15__14_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4971 (
	.O(n3768),
	.A1(n3811),
	.A2(psum2_reg1[15]),
	.B1(n2407),
	.B2(psum2_reg3[15]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4972 (
	.O(n3767),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[15]),
	.C1(n3805),
	.C2(psum4_reg1[15]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4973 (
	.O(n3766),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[15]),
	.C1(n3805),
	.C2(psum3_reg1[15]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U4974 (
	.O(n3765),
	.I1(n3558),
	.I2(psum1_reg3[15]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND4X05AR9 U4975 (
	.O(n3769),
	.I1(n3768),
	.I2(n3767),
	.I3(n3766),
	.I4(n3765), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI12X05AR9 U4976 (
	.O(n3770),
	.A1(n3769),
	.B1(n3802),
	.B2(psum1_reg1[15]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4977 (
	.O(n1489),
	.A1(n3793),
	.A2(n3770),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4978 (
	.O(n1488),
	.A1(n3813),
	.A2(n3770),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4979 (
	.O(n1487),
	.A1(n3814),
	.A2(n3770),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4980 (
	.O(n1486),
	.A1(n3794),
	.A2(n3770),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4981 (
	.O(n1485),
	.A1(n3795),
	.A2(n3770),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4982 (
	.O(n1484),
	.A1(n3817),
	.A2(n3770),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4983 (
	.O(n1483),
	.A1(n2399),
	.A2(n3770),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4984 (
	.O(n1482),
	.A1(n3819),
	.A2(n3770),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4985 (
	.O(n1481),
	.A1(n2400),
	.A2(n3770),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4986 (
	.O(n1480),
	.A1(n3821),
	.A2(n3770),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4987 (
	.O(n1479),
	.A1(n3796),
	.A2(n3770),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4988 (
	.O(n1478),
	.A1(n3797),
	.A2(n3770),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4989 (
	.O(n1477),
	.A1(n3798),
	.A2(n3770),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4990 (
	.O(n1476),
	.A1(n3799),
	.A2(n3770),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4991 (
	.O(n1475),
	.A1(n3825),
	.A2(n3770),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__15_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4992 (
	.O(n1474),
	.A1(n3801),
	.A2(n3770),
	.B1B(Mfifo_psum_M_ffmem_mem_15__15_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4993 (
	.O(n3774),
	.A1(n3811),
	.A2(psum2_reg1[16]),
	.B1(n3751),
	.B2(psum1_reg3[16]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U4994 (
	.O(n3773),
	.A1(n3802),
	.A2(psum1_reg1[16]),
	.B1(n2407),
	.B2(psum2_reg3[16]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4995 (
	.O(n3772),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[16]),
	.C1(n3805),
	.C2(psum3_reg1[16]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U4996 (
	.O(n3771),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[16]),
	.C1(n3805),
	.C2(psum4_reg1[16]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U4997 (
	.O(n3775),
	.I1(n3774),
	.I2(n3773),
	.I3(n3772),
	.I4(n3771), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4998 (
	.O(n1473),
	.A1(n3793),
	.A2(n3775),
	.B1B(n3793),
	.B2B(Mfifo_psum_M_ffmem_mem_0__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U4999 (
	.O(n1472),
	.A1(n3813),
	.A2(n3775),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5000 (
	.O(n1471),
	.A1(n3814),
	.A2(n3775),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5001 (
	.O(n1470),
	.A1(n2398),
	.A2(n3775),
	.B1B(n3794),
	.B2B(Mfifo_psum_M_ffmem_mem_3__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5002 (
	.O(n1469),
	.A1(n3795),
	.A2(n3775),
	.B1B(n3795),
	.B2B(Mfifo_psum_M_ffmem_mem_4__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5003 (
	.O(n1468),
	.A1(n3817),
	.A2(n3775),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5004 (
	.O(n1467),
	.A1(n2399),
	.A2(n3775),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5005 (
	.O(n1466),
	.A1(n3819),
	.A2(n3775),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5006 (
	.O(n1465),
	.A1(n2400),
	.A2(n3775),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5007 (
	.O(n1464),
	.A1(n3821),
	.A2(n3775),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5008 (
	.O(n1463),
	.A1(n3822),
	.A2(n3775),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5009 (
	.O(n1462),
	.A1(n3797),
	.A2(n3775),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5010 (
	.O(n1461),
	.A1(n3798),
	.A2(n3775),
	.B1B(n3798),
	.B2B(Mfifo_psum_M_ffmem_mem_12__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5011 (
	.O(n1460),
	.A1(n3799),
	.A2(n3775),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5012 (
	.O(n1459),
	.A1(n3825),
	.A2(n3775),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__16_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5013 (
	.O(n1458),
	.A1(n3801),
	.A2(n3775),
	.B1B(Mfifo_psum_M_ffmem_mem_15__16_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   LOWMUX2X05AR9 U5014 (
	.O(n3782),
	.EB(n3776),
	.I0(psum4_reg3[17]),
	.I1(psum4_reg1[17]),
	.S(sel_ccp), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   INVX05AR9 U5015 (
	.O(n3779),
	.I(psum2_reg1[17]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U5016 (
	.O(n3778),
	.A1(n3751),
	.A2(psum1_reg3[17]),
	.B1(n3802),
	.B2(psum1_reg1[17]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U5017 (
	.O(n3777),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[17]),
	.C1(n3805),
	.C2(psum3_reg1[17]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI112X05AR9 U5018 (
	.O(n3781),
	.A1(n3778),
	.B1(n3777),
	.C1(n3780),
	.C2(n3779), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5019 (
	.O(n1457),
	.A1(n3793),
	.A2(n3783),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5020 (
	.O(n1456),
	.A1(n3813),
	.A2(n3783),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5021 (
	.O(n1455),
	.A1(n3814),
	.A2(n3783),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5022 (
	.O(n1454),
	.A1(n3794),
	.A2(n3783),
	.B1B(n3794),
	.B2B(Mfifo_psum_M_ffmem_mem_3__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5023 (
	.O(n1453),
	.A1(n3795),
	.A2(n3783),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5024 (
	.O(n1452),
	.A1(n3817),
	.A2(n3783),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5025 (
	.O(n1451),
	.A1(n2399),
	.A2(n3783),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5026 (
	.O(n1450),
	.A1(n3819),
	.A2(n3783),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5027 (
	.O(n1449),
	.A1(n2400),
	.A2(n3783),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5028 (
	.O(n1448),
	.A1(n3821),
	.A2(n3783),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5029 (
	.O(n1447),
	.A1(n3796),
	.A2(n3783),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5030 (
	.O(n1446),
	.A1(n3797),
	.A2(n3783),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5031 (
	.O(n1445),
	.A1(n3798),
	.A2(n3783),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5032 (
	.O(n1444),
	.A1(n3799),
	.A2(n3783),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5033 (
	.O(n1443),
	.A1(n3825),
	.A2(n3783),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__17_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5034 (
	.O(n1442),
	.A1(n3801),
	.A2(n3783),
	.B1B(Mfifo_psum_M_ffmem_mem_15__17_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U5035 (
	.O(n3787),
	.A1(n3811),
	.A2(psum2_reg1[18]),
	.B1(n3802),
	.B2(psum1_reg1[18]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U5036 (
	.O(n3786),
	.A1(n3558),
	.A2(psum1_reg3[18]),
	.B1(n2407),
	.B2(psum2_reg3[18]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U5037 (
	.O(n3785),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[18]),
	.C1(n3805),
	.C2(psum4_reg1[18]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U5038 (
	.O(n3784),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[18]),
	.C1(n3805),
	.C2(psum3_reg1[18]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U5039 (
	.O(n3788),
	.I1(n3787),
	.I2(n3786),
	.I3(n3785),
	.I4(n3784), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5040 (
	.O(n1441),
	.A1(n3793),
	.A2(n3788),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5041 (
	.O(n1440),
	.A1(n3813),
	.A2(n3788),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5042 (
	.O(n1439),
	.A1(n3814),
	.A2(n3788),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5043 (
	.O(n1438),
	.A1(n2398),
	.A2(n3788),
	.B1B(n3794),
	.B2B(Mfifo_psum_M_ffmem_mem_3__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5044 (
	.O(n1437),
	.A1(n3795),
	.A2(n3788),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5045 (
	.O(n1436),
	.A1(n3817),
	.A2(n3788),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5046 (
	.O(n1435),
	.A1(n2399),
	.A2(n3788),
	.B1B(n3818),
	.B2B(Mfifo_psum_M_ffmem_mem_6__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5047 (
	.O(n1434),
	.A1(n3819),
	.A2(n3788),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5048 (
	.O(n1433),
	.A1(n2400),
	.A2(n3788),
	.B1B(n3820),
	.B2B(Mfifo_psum_M_ffmem_mem_8__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5049 (
	.O(n1432),
	.A1(n3821),
	.A2(n3788),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5050 (
	.O(n1431),
	.A1(n3822),
	.A2(n3788),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5051 (
	.O(n1430),
	.A1(n3797),
	.A2(n3788),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5052 (
	.O(n1429),
	.A1(n3798),
	.A2(n3788),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5053 (
	.O(n1428),
	.A1(n3799),
	.A2(n3788),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5054 (
	.O(n1427),
	.A1(n3825),
	.A2(n3788),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__18_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5055 (
	.O(n1426),
	.A1(n3801),
	.A2(n3788),
	.B1B(Mfifo_psum_M_ffmem_mem_15__18_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U5056 (
	.O(n3792),
	.A1(n3558),
	.A2(psum1_reg3[19]),
	.B1(n3802),
	.B2(psum1_reg1[19]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U5057 (
	.O(n3791),
	.A1(n3811),
	.A2(psum2_reg1[19]),
	.B1(n2407),
	.B2(psum2_reg3[19]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U5058 (
	.O(n3790),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[19]),
	.C1(n3805),
	.C2(psum4_reg1[19]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U5059 (
	.O(n3789),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[19]),
	.C1(n3805),
	.C2(psum3_reg1[19]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AND4X05AR9 U5060 (
	.O(n3800),
	.I1(n3792),
	.I2(n3791),
	.I3(n3790),
	.I4(n3789), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5061 (
	.O(n1425),
	.A1(n3793),
	.A2(n3800),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5062 (
	.O(n1424),
	.A1(n3813),
	.A2(n3800),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5063 (
	.O(n1423),
	.A1(n3814),
	.A2(n3800),
	.B1B(n3815),
	.B2B(Mfifo_psum_M_ffmem_mem_2__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5064 (
	.O(n1422),
	.A1(n2398),
	.A2(n3800),
	.B1B(n3794),
	.B2B(Mfifo_psum_M_ffmem_mem_3__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5065 (
	.O(n1421),
	.A1(n3795),
	.A2(n3800),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5066 (
	.O(n1420),
	.A1(n3817),
	.A2(n3800),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5067 (
	.O(n1419),
	.A1(n2399),
	.A2(n3800),
	.B1B(n3818),
	.B2B(Mfifo_psum_M_ffmem_mem_6__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5068 (
	.O(n1418),
	.A1(n3819),
	.A2(n3800),
	.B1B(n3819),
	.B2B(Mfifo_psum_M_ffmem_mem_7__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5069 (
	.O(n1417),
	.A1(n2400),
	.A2(n3800),
	.B1B(n3820),
	.B2B(Mfifo_psum_M_ffmem_mem_8__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5070 (
	.O(n1416),
	.A1(n3821),
	.A2(n3800),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5071 (
	.O(n1415),
	.A1(n3822),
	.A2(n3800),
	.B1B(n3796),
	.B2B(Mfifo_psum_M_ffmem_mem_10__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5072 (
	.O(n1414),
	.A1(n3797),
	.A2(n3800),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5073 (
	.O(n1413),
	.A1(n3798),
	.A2(n3800),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5074 (
	.O(n1412),
	.A1(n3799),
	.A2(n3800),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5075 (
	.O(n1411),
	.A1(n3824),
	.A2(n3800),
	.B1B(n3825),
	.B2B(Mfifo_psum_M_ffmem_mem_14__19_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5076 (
	.O(n1410),
	.A1(n3801),
	.A2(n3800),
	.B1B(Mfifo_psum_M_ffmem_mem_15__19_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22X05AR9 U5077 (
	.O(n3809),
	.A1(n3802),
	.A2(psum1_reg1[20]),
	.B1(n2407),
	.B2(psum2_reg3[20]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U5078 (
	.O(n3808),
	.A1(n3803),
	.B1(sel_ccp),
	.B2(psum3_reg3[20]),
	.C1(n3805),
	.C2(psum3_reg1[20]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI122X05AR9 U5079 (
	.O(n3807),
	.A1(n3640),
	.B1(sel_ccp),
	.B2(psum4_reg3[20]),
	.C1(n3805),
	.C2(psum4_reg1[20]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U5080 (
	.O(n3806),
	.I1(n3558),
	.I2(psum1_reg3[20]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5081 (
	.O(n1409),
	.A1(n3812),
	.A2(n3826),
	.B1B(n3812),
	.B2B(Mfifo_psum_M_ffmem_mem_0__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5082 (
	.O(n1408),
	.A1(n3813),
	.A2(n3826),
	.B1B(n3813),
	.B2B(Mfifo_psum_M_ffmem_mem_1__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5083 (
	.O(n1407),
	.A1(n3815),
	.A2(n3826),
	.B1B(n3814),
	.B2B(Mfifo_psum_M_ffmem_mem_2__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5084 (
	.O(n1406),
	.A1(n2398),
	.A2(n3826),
	.B1B(n2398),
	.B2B(Mfifo_psum_M_ffmem_mem_3__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5085 (
	.O(n1405),
	.A1(n3816),
	.A2(n3826),
	.B1B(n3816),
	.B2B(Mfifo_psum_M_ffmem_mem_4__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5086 (
	.O(n1404),
	.A1(n3817),
	.A2(n3826),
	.B1B(n3817),
	.B2B(Mfifo_psum_M_ffmem_mem_5__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5087 (
	.O(n1403),
	.A1(n3818),
	.A2(n3826),
	.B1B(n2399),
	.B2B(Mfifo_psum_M_ffmem_mem_6__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5088 (
	.O(n1402),
	.A1(n3819),
	.A2(n3826),
	.B1B(n3738),
	.B2B(Mfifo_psum_M_ffmem_mem_7__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5089 (
	.O(n1401),
	.A1(n3820),
	.A2(n3826),
	.B1B(n2400),
	.B2B(Mfifo_psum_M_ffmem_mem_8__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5090 (
	.O(n1400),
	.A1(n3821),
	.A2(n3826),
	.B1B(n3821),
	.B2B(Mfifo_psum_M_ffmem_mem_9__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5091 (
	.O(n1399),
	.A1(n3822),
	.A2(n3826),
	.B1B(n3822),
	.B2B(Mfifo_psum_M_ffmem_mem_10__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5092 (
	.O(n1398),
	.A1(n3797),
	.A2(n3826),
	.B1B(n3797),
	.B2B(Mfifo_psum_M_ffmem_mem_11__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5093 (
	.O(n1397),
	.A1(n3823),
	.A2(n3826),
	.B1B(n3823),
	.B2B(Mfifo_psum_M_ffmem_mem_12__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5094 (
	.O(n1396),
	.A1(n3799),
	.A2(n3826),
	.B1B(n3799),
	.B2B(Mfifo_psum_M_ffmem_mem_13__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5095 (
	.O(n1395),
	.A1(n3825),
	.A2(n3826),
	.B1B(n3824),
	.B2B(Mfifo_psum_M_ffmem_mem_14__20_), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   AOI22B2X05AR9 U5096 (
	.O(n1394),
	.A1(n3801),
	.A2(n3826),
	.B1B(Mfifo_psum_M_ffmem_mem_15__20_),
	.B2B(n3801), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   NAND2X05AR9 U5097 (
	.O(n3828),
	.I1(n3827),
	.I2(int_kx[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));
   OAI12B2X05AR9 U5098 (
	.O(n1393),
	.A1(n3828),
	.B1B(n3829),
	.B2B(Mcntl_Mcntldata_kx_reg[1]), 
	.VCCK(VCCK), 
	.GNDK(GNDK));

   // Fillers and physical instances.
   FILLERC16CR9 ENDCAP_948 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_947 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_946 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_945 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_944 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_943 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_942 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_941 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_940 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_939 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_938 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_937 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_936 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_935 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_934 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_933 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_932 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_931 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_930 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_929 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_928 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_927 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_926 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_925 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_924 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_923 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_922 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_921 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_920 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_919 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_918 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_917 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_916 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_915 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_914 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_913 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_912 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_911 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_910 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_909 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_908 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_907 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_906 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_905 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_904 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_903 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_902 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_901 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_900 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_899 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_898 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_897 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_896 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_895 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_894 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_893 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_892 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_891 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_890 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_889 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_888 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_887 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_886 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_885 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_884 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_883 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_882 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_881 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_880 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_879 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_878 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_877 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_876 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_875 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_874 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_873 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_872 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_871 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_870 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_869 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_868 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_867 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_866 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_865 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_864 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_863 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_862 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_861 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_860 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_859 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_858 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_857 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_856 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_855 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_854 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_853 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_852 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_851 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_850 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_849 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_848 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_847 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_846 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_845 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_844 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_843 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_842 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_841 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_840 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_839 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_838 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_837 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_836 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_835 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_834 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_833 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_832 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_831 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_830 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_829 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_828 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_827 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_826 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_825 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_824 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_823 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_822 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_821 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_820 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_819 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_818 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_817 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_816 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_815 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_814 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_813 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_812 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_811 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_810 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_809 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_808 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_807 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_806 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_805 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_804 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_803 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_802 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_801 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_800 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_799 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_798 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_797 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_796 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_795 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_794 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_793 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_792 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_791 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_790 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_789 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_788 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_787 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_786 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_785 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_784 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_783 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_782 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_781 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_780 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_779 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_778 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_777 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_776 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_775 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_774 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_773 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_772 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_771 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_770 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_769 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_768 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_767 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_766 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_765 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_764 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_763 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_762 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_761 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_760 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_759 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_758 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_757 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_756 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_755 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_754 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_753 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_752 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_751 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_750 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_749 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_748 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_747 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_746 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_745 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_744 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_743 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_742 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_741 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_740 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_739 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_738 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_737 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_736 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_735 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_734 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_733 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_732 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_731 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_730 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_729 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_728 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_727 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_726 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_725 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_724 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_723 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_722 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_721 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_720 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_719 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_718 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_717 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_716 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_715 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_714 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_713 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_712 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_711 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_710 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_709 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_708 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_707 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_706 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_705 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_704 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_703 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_702 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_701 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_700 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_699 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_698 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_697 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_696 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_695 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_694 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_693 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_692 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_691 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_690 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_689 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_688 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_687 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_686 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_685 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_684 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_683 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_682 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_681 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_680 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_679 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_678 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_677 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_676 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_675 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_674 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_673 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_672 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_671 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_670 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_669 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_668 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_667 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_666 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_665 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_664 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_663 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_662 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_661 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_660 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_659 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_658 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_657 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_656 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_655 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_654 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_653 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_652 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_651 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_650 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_649 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_648 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_647 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_646 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_645 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_644 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_643 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_642 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_641 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_640 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_639 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_638 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_637 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_636 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_635 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_634 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_633 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_632 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_631 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_630 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_629 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_628 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_627 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_626 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_625 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_624 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_623 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_622 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_621 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_620 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_619 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_618 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_617 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_616 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_615 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_614 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_613 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_612 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_611 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_610 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_609 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_608 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_607 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_606 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_605 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_604 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_603 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_602 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_601 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_600 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_599 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_598 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_597 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_596 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_595 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_594 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_593 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_592 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_591 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_590 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_589 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_588 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_587 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_586 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_585 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_584 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_583 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_582 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_581 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_580 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_579 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_578 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_577 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_576 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_575 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_574 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_573 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_572 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_571 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_570 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_569 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_568 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_567 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_566 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_565 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_564 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_563 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_562 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_561 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_560 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_559 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_558 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_557 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_556 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_555 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_554 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_553 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_552 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_551 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_550 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_549 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_548 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_547 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_546 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_545 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_544 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_543 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_542 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_541 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_540 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_539 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_538 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_537 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_536 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_535 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_534 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_533 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_532 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_531 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_530 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_529 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_528 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_527 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_526 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_525 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_524 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_523 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_522 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_521 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_520 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_519 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_518 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_517 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_516 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_515 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_514 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_513 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_512 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_511 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_510 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_509 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_508 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_507 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_506 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_505 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_504 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_503 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_502 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_501 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_500 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_499 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_498 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_497 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_496 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_495 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_494 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_493 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_492 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_491 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_490 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_489 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_488 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_487 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_486 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_485 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_484 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_483 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_482 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_481 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_480 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_479 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_478 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_477 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_476 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_475 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_474 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_473 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_472 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_471 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_470 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_469 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_468 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_467 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_466 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_465 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_464 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_463 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_462 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_461 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_460 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_459 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_458 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_457 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_456 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_455 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_454 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_453 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_452 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_451 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_450 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_449 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_448 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_447 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_446 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_445 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_444 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_443 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_442 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_441 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_440 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_439 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_438 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_437 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_436 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_435 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_434 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_433 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_432 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_431 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_430 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_429 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_428 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_427 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_426 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_425 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_424 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_423 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_422 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_421 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_420 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_419 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_418 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_417 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_416 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_415 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_414 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_413 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_412 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_411 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_410 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_409 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_408 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_407 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_406 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_405 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_404 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_403 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_402 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_401 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_400 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_399 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_398 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_397 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_396 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_395 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_394 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_393 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_392 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_391 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_390 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_389 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_388 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_387 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_386 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_385 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_384 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_383 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_382 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_381 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_380 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_379 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_378 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_377 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_376 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_375 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_374 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_373 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_372 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_371 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_370 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_369 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_368 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_367 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_366 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_365 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_364 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_363 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_362 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_361 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_360 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_359 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_358 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_357 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_356 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_355 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_354 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_353 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_352 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_351 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_350 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_349 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_348 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_347 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_346 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_345 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_344 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_343 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_342 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_341 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_340 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_339 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_338 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_337 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_336 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_335 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_334 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_333 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_332 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_331 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_330 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_329 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_328 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_327 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_326 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_325 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_324 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_323 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_322 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_321 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_320 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_319 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_318 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_317 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_316 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_315 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_314 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_313 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_312 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_311 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_310 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_309 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_308 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_307 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_306 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_305 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_304 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_303 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_302 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_301 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_300 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_299 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_298 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_297 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_296 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_295 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_294 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_293 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_292 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_291 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_290 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_289 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_288 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_287 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_286 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_285 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_284 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_283 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_282 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_281 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_280 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_279 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_278 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_277 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_276 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_275 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_274 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_273 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_272 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_271 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_270 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_269 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_268 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_267 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_266 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_265 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_264 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_263 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_262 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_261 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_260 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_259 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_258 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_257 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_256 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_255 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_254 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_253 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_252 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_251 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_250 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_249 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_248 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_247 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_246 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_245 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_244 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_243 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_242 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_241 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_240 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_239 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_238 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_237 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_236 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_235 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_234 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_233 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_232 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_231 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_230 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_229 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_228 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_227 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_226 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_225 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_224 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_223 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_222 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_221 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_220 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_219 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_218 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_217 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_216 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_215 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_214 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_213 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_212 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_211 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_210 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_209 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_208 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_207 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_206 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_205 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_204 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_203 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_202 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_201 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_200 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_199 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_198 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_197 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_196 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_195 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_194 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_193 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_192 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_191 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_190 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_189 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_188 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_187 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_186 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_185 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_184 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_183 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_182 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_181 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_180 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_179 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_178 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_177 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_176 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_175 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_174 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_173 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_172 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_171 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_170 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_169 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_168 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_167 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_166 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_165 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_164 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_163 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_162 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_161 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_160 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_159 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_158 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_157 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_156 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_155 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_154 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_153 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_152 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_151 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_150 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_149 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_148 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_147 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_146 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_145 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_144 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_143 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_142 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_141 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_140 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_139 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_138 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_137 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_136 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_135 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_134 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_133 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_132 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_131 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_130 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_129 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_128 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_127 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_126 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_125 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_124 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_123 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_122 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_121 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_120 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_119 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_118 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_117 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_116 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_115 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_114 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_113 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_112 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_111 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_110 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_109 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_108 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_107 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_106 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_105 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_104 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_103 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_102 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_101 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_100 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_99 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_98 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_97 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_96 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_95 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_94 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_93 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_92 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_91 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_90 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_89 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_88 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_87 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_86 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_85 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_84 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_83 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_82 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_81 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_80 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_79 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_78 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_77 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_76 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_75 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_74 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_73 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_72 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_71 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_70 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_69 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_68 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_67 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_66 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_65 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_64 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_63 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_62 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_61 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_60 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_59 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_58 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_57 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_56 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_55 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_54 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_53 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_52 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_51 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_50 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_49 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_48 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_47 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_46 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_45 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_44 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_43 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_42 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_41 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_40 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_39 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_38 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_37 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_36 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_35 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_34 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_33 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_32 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_31 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_30 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_29 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_28 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_27 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_26 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_25 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_24 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_23 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_22 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_21 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_20 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_19 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_18 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_17 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_16 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_15 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_14 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_13 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_12 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_11 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_10 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_9 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_8 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_7 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_6 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_5 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_4 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_3 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_2 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
   FILLERC16CR9 ENDCAP_1 (
	.VCCK(VCCK), 
	.GNDK(GNDK) );
endmodule
